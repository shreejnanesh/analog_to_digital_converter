
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41_USR1.7.43
#
# TECH LIB NAME: gsclib090
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 2000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
## Site is specified in gsclib090 tech file; and there is no need here.
## Make sure to correct the "SITE" value to 'gsclib090site' on each macro cell.
#SITE gsclib090site
#    SYMMETRY Y  ;
#    CLASS core  ;
#    SIZE 0.2900 BY 2.6100 ;
#END gsclib090site

MACRO XOR3XL
    CLASS CORE ;
    FOREIGN XOR3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3684  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2700 1.5600 8.5100 2.2500 ;
        RECT  8.3900 0.3600 8.5100 2.2500 ;
        RECT  8.1350 0.6500 8.5100 0.8000 ;
        RECT  8.2700 0.3600 8.5100 0.8000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0840  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.0700 0.3250 1.4700 ;
        RECT  0.0700 1.1750 0.3250 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3168  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2520  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.2571  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        RECT  0.8450 1.0300 1.0250 1.3750 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0800 1.3500 6.8100 1.4700 ;
        RECT  6.0800 1.2300 6.3650 1.4700 ;
        RECT  6.0800 0.9050 6.2000 1.4700 ;
        RECT  5.6950 0.9050 6.2000 1.0250 ;
        END
    END C
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.7300 2.2900 7.9700 2.7900 ;
        RECT  7.7900 1.6900 7.9100 2.7900 ;
        RECT  1.8650 2.2700 2.1050 2.7900 ;
        RECT  0.6850 2.2900 0.9250 2.7900 ;
        RECT  0.7450 1.9700 0.8650 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.7300 -0.1800 7.9700 0.3200 ;
        RECT  7.7900 -0.1800 7.9100 0.6700 ;
        RECT  1.8650 -0.1800 2.1050 0.3200 ;
        RECT  0.6850 -0.1800 0.9250 0.3200 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  8.2300 1.3150 7.6700 1.3150 7.6700 2.1700 6.2600 2.1700 6.2600 1.8900 6.5600 1.8900
                 6.5600 2.0500 7.5500 2.0500 7.5500 0.6200 7.4200 0.6200 7.4200 0.4800 6.2600 0.4800
                 6.2600 0.3600 7.5400 0.3600 7.5400 0.5000 7.6700 0.5000 7.6700 1.1950 7.9900 1.1950
                 7.9900 1.0750 8.2300 1.0750 ;
        POLYGON  7.4300 0.8600 7.3450 0.8600 7.3450 1.8100 7.4300 1.8100 7.4300 1.9300 7.1900 1.9300
                 7.1900 1.8100 7.2250 1.8100 7.2250 0.8600 7.1900 0.8600 7.1900 0.7400 7.4300 0.7400 ;
        POLYGON  7.0500 1.7700 7.0400 1.7700 7.0400 1.7900 6.8000 1.7900 6.8000 1.7700 4.2750 1.7700
                 4.2750 1.6500 5.0950 1.6500 5.0950 0.7200 4.2700 0.7200 4.2700 0.6000 5.2150 0.6000
                 5.2150 1.6500 6.9300 1.6500 6.9300 0.7200 6.8000 0.7200 6.8000 0.6000 7.0500 0.6000 ;
        POLYGON  5.9600 0.7050 5.9000 0.7050 5.9000 0.7200 5.4800 0.7200 5.4800 1.4050 5.9600 1.4050
                 5.9600 1.5250 5.3600 1.5250 5.3600 0.6000 5.7200 0.6000 5.7200 0.5850 5.9600 0.5850 ;
        RECT  2.9850 1.8900 5.9600 2.0100 ;
        RECT  2.4050 0.3600 5.6400 0.4800 ;
        RECT  2.4050 2.1300 5.6400 2.2500 ;
        POLYGON  4.8400 1.0400 4.1700 1.0400 4.1700 1.4150 4.0500 1.4150 4.0500 0.9200 4.8400 0.9200 ;
        POLYGON  3.9850 0.7200 3.8400 0.7200 3.8400 1.7700 1.7250 1.7700 1.7250 2.1700 0.9850 2.1700
                 0.9850 1.8100 0.3250 1.8100 0.3250 1.9300 0.1450 1.9300 0.1450 1.6900 0.5050 1.6900
                 0.5050 0.9200 0.2050 0.9200 0.2050 0.4400 1.6050 0.4400 1.6050 0.3200 1.7250 0.3200
                 1.7250 0.5600 0.3250 0.5600 0.3250 0.8000 0.6250 0.8000 0.6250 1.6900 1.1050 1.6900
                 1.1050 2.0500 1.6050 2.0500 1.6050 1.6500 3.7200 1.6500 3.7200 0.6000 3.9850 0.6000 ;
        POLYGON  3.5850 1.0400 3.4050 1.0400 3.4050 1.0000 2.8100 1.0000 2.8100 1.1600 2.8850 1.1600
                 2.8850 1.2800 2.6450 1.2800 2.6450 1.1600 2.6900 1.1600 2.6900 0.8800 3.4050 0.8800
                 3.4050 0.8000 3.5850 0.8000 ;
        POLYGON  3.2250 1.5300 1.9400 1.5300 1.9400 0.6000 3.2050 0.6000 3.2050 0.7200 2.0600 0.7200
                 2.0600 1.4100 3.2250 1.4100 ;
        POLYGON  1.4850 1.1200 1.4050 1.1200 1.4050 1.8100 1.4650 1.8100 1.4650 1.9300 1.2250 1.9300
                 1.2250 1.8100 1.2850 1.8100 1.2850 1.1200 1.2450 1.1200 1.2450 1.0000 1.2850 1.0000
                 1.2850 0.8000 1.2250 0.8000 1.2250 0.6800 1.4650 0.6800 1.4650 0.8000 1.4050 0.8000
                 1.4050 1.0000 1.4850 1.0000 ;
    END
END XOR3XL

MACRO XOR3X1
    CLASS CORE ;
    FOREIGN XOR3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4014  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2700 1.5600 8.5100 2.2500 ;
        RECT  8.3900 0.3600 8.5100 2.2500 ;
        RECT  8.1350 0.6500 8.5100 0.8000 ;
        RECT  8.2700 0.3600 8.5100 0.8000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0990  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.0700 0.3250 1.4700 ;
        RECT  0.0700 1.1750 0.3250 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3198  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2670  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.1978  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        RECT  0.8450 1.0300 1.0250 1.3750 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0800 1.3500 6.8100 1.4700 ;
        RECT  6.0800 1.2300 6.3650 1.4700 ;
        RECT  6.0800 0.9050 6.2000 1.4700 ;
        RECT  5.6950 0.9050 6.2000 1.0250 ;
        END
    END C
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.7300 2.2900 7.9700 2.7900 ;
        RECT  7.7900 1.6900 7.9100 2.7900 ;
        RECT  1.8650 2.2700 2.1050 2.7900 ;
        RECT  0.6850 2.2900 0.9250 2.7900 ;
        RECT  0.7450 1.9700 0.8650 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.7300 -0.1800 7.9700 0.3200 ;
        RECT  7.7900 -0.1800 7.9100 0.6700 ;
        RECT  1.8650 -0.1800 2.1050 0.3200 ;
        RECT  0.6850 -0.1800 0.9250 0.3200 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  8.2300 1.3150 7.6700 1.3150 7.6700 2.1700 6.2600 2.1700 6.2600 1.8900 6.5600 1.8900
                 6.5600 2.0500 7.5500 2.0500 7.5500 0.6200 7.4200 0.6200 7.4200 0.4800 6.2600 0.4800
                 6.2600 0.3600 7.5400 0.3600 7.5400 0.5000 7.6700 0.5000 7.6700 1.1950 7.9900 1.1950
                 7.9900 1.0750 8.2300 1.0750 ;
        POLYGON  7.4300 0.8600 7.3450 0.8600 7.3450 1.8100 7.4300 1.8100 7.4300 1.9300 7.1900 1.9300
                 7.1900 1.8100 7.2250 1.8100 7.2250 0.8600 7.1900 0.8600 7.1900 0.7400 7.4300 0.7400 ;
        POLYGON  7.0500 1.7700 7.0400 1.7700 7.0400 1.7900 6.8000 1.7900 6.8000 1.7700 4.2750 1.7700
                 4.2750 1.6500 5.0950 1.6500 5.0950 0.7200 4.5250 0.7200 4.5250 0.6000 5.2150 0.6000
                 5.2150 1.6500 6.9300 1.6500 6.9300 0.7200 6.8000 0.7200 6.8000 0.6000 7.0500 0.6000 ;
        POLYGON  5.9600 0.7050 5.9000 0.7050 5.9000 0.7200 5.4800 0.7200 5.4800 1.4050 5.9600 1.4050
                 5.9600 1.5250 5.3600 1.5250 5.3600 0.6000 5.7200 0.6000 5.7200 0.5850 5.9600 0.5850 ;
        RECT  2.9850 1.8900 5.9600 2.0100 ;
        RECT  2.4050 0.3600 5.6400 0.4800 ;
        RECT  2.4050 2.1300 5.6400 2.2500 ;
        POLYGON  4.9700 1.0400 4.1700 1.0400 4.1700 1.2850 4.0500 1.2850 4.0500 0.9200 4.9700 0.9200 ;
        POLYGON  4.0750 0.7200 3.9300 0.7200 3.9300 1.7700 1.7250 1.7700 1.7250 2.1700 0.9850 2.1700
                 0.9850 1.8100 0.3250 1.8100 0.3250 1.9300 0.2050 1.9300 0.2050 1.6900 0.5050 1.6900
                 0.5050 0.9200 0.2050 0.9200 0.2050 0.4400 1.6050 0.4400 1.6050 0.3200 1.7250 0.3200
                 1.7250 0.5600 0.3250 0.5600 0.3250 0.8000 0.6250 0.8000 0.6250 1.6900 1.1050 1.6900
                 1.1050 2.0500 1.6050 2.0500 1.6050 1.6500 3.8100 1.6500 3.8100 0.6000 4.0750 0.6000 ;
        POLYGON  3.6900 1.0800 3.5700 1.0800 3.5700 1.0200 2.8100 1.0200 2.8100 1.1600 2.8850 1.1600
                 2.8850 1.2800 2.6450 1.2800 2.6450 1.1600 2.6900 1.1600 2.6900 0.9000 3.5700 0.9000
                 3.5700 0.8400 3.6900 0.8400 ;
        POLYGON  3.2250 1.5300 1.9400 1.5300 1.9400 0.6000 3.2050 0.6000 3.2050 0.7200 2.0600 0.7200
                 2.0600 1.4100 3.2250 1.4100 ;
        POLYGON  1.4850 1.1200 1.4050 1.1200 1.4050 1.8100 1.4650 1.8100 1.4650 1.9300 1.2250 1.9300
                 1.2250 1.8100 1.2850 1.8100 1.2850 1.1200 1.2450 1.1200 1.2450 1.0000 1.2850 1.0000
                 1.2850 0.8000 1.2250 0.8000 1.2250 0.6800 1.4650 0.6800 1.4650 0.8000 1.4050 0.8000
                 1.4050 1.0000 1.4850 1.0000 ;
    END
END XOR3X1

MACRO XOR2XL
    CLASS CORE ;
    FOREIGN XOR2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8350 1.2900 0.9550 1.5300 ;
        RECT  0.6800 1.4100 0.9550 1.5300 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4150 1.2700 2.6550 1.3900 ;
        RECT  1.3350 1.1700 2.5350 1.2900 ;
        RECT  1.8550 1.0900 2.0950 1.2900 ;
        RECT  1.7550 1.1700 2.0150 1.3800 ;
        RECT  1.3350 1.1700 1.4550 1.5500 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.5500 0.2550 1.8700 ;
        RECT  0.0700 1.4650 0.2550 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.3550 0.6100 2.5950 0.7300 ;
        RECT  2.3550 -0.1800 2.4750 0.7300 ;
        RECT  0.4950 0.6100 0.7350 0.7300 ;
        RECT  0.4950 -0.1800 0.6150 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.2150 1.7500 2.3350 2.7900 ;
        RECT  0.6150 2.2300 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.9550 0.7900 2.8950 0.7900 2.8950 1.7500 2.7550 1.7500 2.7550 1.8700 2.6350 1.8700
                 2.6350 1.6300 1.8950 1.6300 1.8950 2.2500 1.6550 2.2500 1.6550 2.1300 1.7750 2.1300
                 1.7750 1.5100 2.7750 1.5100 2.7750 0.6700 2.8350 0.6700 2.8350 0.5500 2.9550 0.5500 ;
        POLYGON  2.4550 1.0500 2.2150 1.0500 2.2150 0.9700 1.2150 0.9700 1.2150 1.8700 1.0950 1.8700
                 1.0950 0.6100 1.3350 0.6100 1.3350 0.7300 1.2150 0.7300 1.2150 0.8500 2.3350 0.8500
                 2.3350 0.9300 2.4550 0.9300 ;
        POLYGON  1.9550 0.7300 1.7150 0.7300 1.7150 0.4900 0.9750 0.4900 0.9750 1.1700 0.5300 1.1700
                 0.5300 1.8450 0.7400 1.8450 0.7400 1.9900 1.4150 1.9900 1.4150 1.8700 1.5150 1.8700
                 1.5150 1.7500 1.6350 1.7500 1.6350 1.9900 1.5350 1.9900 1.5350 2.1100 0.6200 2.1100
                 0.6200 1.9650 0.4100 1.9650 0.4100 0.9500 0.5300 0.9500 0.5300 1.0500 0.8550 1.0500
                 0.8550 0.3700 1.8350 0.3700 1.8350 0.6100 1.9550 0.6100 ;
    END
END XOR2XL

MACRO XOR2X4
    CLASS CORE ;
    FOREIGN XOR2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.1800 2.1750 1.3450 ;
        RECT  1.7550 1.1800 2.0150 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7950 0.9400 3.9150 1.1800 ;
        RECT  3.0150 0.9700 3.9150 1.0900 ;
        RECT  3.4950 0.9400 3.9150 1.0900 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 1.7400 1.5750 2.2100 ;
        RECT  1.2150 0.7000 1.5150 0.8200 ;
        RECT  1.3950 0.5800 1.5150 0.8200 ;
        RECT  1.2750 1.7400 1.5750 1.8600 ;
        RECT  1.2750 1.3200 1.3950 1.8600 ;
        RECT  0.6500 0.8400 1.3350 0.9600 ;
        RECT  1.2150 0.7000 1.3350 0.9600 ;
        RECT  0.6500 1.3200 1.3950 1.4400 ;
        RECT  0.6500 1.1750 0.8000 1.4400 ;
        RECT  0.6500 0.7300 0.7700 1.5600 ;
        RECT  0.6150 1.4400 0.7350 2.2100 ;
        RECT  0.4950 0.7300 0.7700 0.8500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.5350 0.4600 3.7750 0.5800 ;
        RECT  3.5350 -0.1800 3.6550 0.5800 ;
        RECT  1.8150 -0.1800 1.9350 0.7200 ;
        RECT  0.9750 -0.1800 1.0950 0.7200 ;
        RECT  0.1350 -0.1800 0.2550 0.7200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.5950 1.7700 3.7150 2.7900 ;
        RECT  1.8150 2.0100 2.0550 2.1500 ;
        RECT  1.8150 2.0100 1.9350 2.7900 ;
        RECT  1.0350 1.5600 1.1550 2.7900 ;
        RECT  0.1950 1.5600 0.3150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.1550 1.8900 4.1350 1.8900 4.1350 2.0100 4.0150 2.0100 4.0150 1.7700 4.0350 1.7700
                 4.0350 0.8200 2.8950 0.8200 2.8950 1.2900 3.2750 1.2900 3.2750 1.4100 2.7750 1.4100
                 2.7750 1.0500 2.6550 1.0500 2.6550 1.1700 2.5350 1.1700 2.5350 0.9300 2.7750 0.9300
                 2.7750 0.7000 4.0150 0.7000 4.0150 0.4000 4.1350 0.4000 4.1350 0.5200 4.1550 0.5200 ;
        POLYGON  3.6350 1.4100 3.5150 1.4100 3.5150 1.6500 2.6550 1.6500 2.6550 2.0100 2.5350 2.0100
                 2.5350 1.6500 2.2950 1.6500 2.2950 0.6500 2.5550 0.6500 2.5550 0.7700 2.4150 0.7700
                 2.4150 1.5300 3.3950 1.5300 3.3950 1.2900 3.6350 1.2900 ;
        POLYGON  3.0750 2.2500 2.1750 2.2500 2.1750 1.8900 1.9100 1.8900 1.9100 1.6200 1.5150 1.6200
                 1.5150 1.2000 1.2550 1.2000 1.2550 1.0800 1.5150 1.0800 1.5150 0.9400 2.0550 0.9400
                 2.0550 0.4100 2.8550 0.4100 2.8550 0.4600 2.9750 0.4600 2.9750 0.5800 2.7350 0.5800
                 2.7350 0.5300 2.1750 0.5300 2.1750 1.0600 1.6350 1.0600 1.6350 1.5000 2.0300 1.5000
                 2.0300 1.7700 2.2950 1.7700 2.2950 2.1300 2.9550 2.1300 2.9550 1.7700 3.0750 1.7700 ;
    END
END XOR2X4

MACRO XOR2X2
    CLASS CORE ;
    FOREIGN XOR2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 1.2200 1.3350 1.4600 ;
        RECT  0.8850 1.2300 1.3350 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8150 1.1800 3.1750 1.3000 ;
        RECT  2.3350 1.1800 2.5950 1.3800 ;
        RECT  2.2550 1.1400 2.4950 1.3000 ;
        RECT  1.6950 1.3400 1.9350 1.4600 ;
        RECT  1.8150 1.1800 1.9350 1.4600 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.7400 0.7150 2.2100 ;
        RECT  0.4050 0.7400 0.6750 0.8600 ;
        RECT  0.5550 0.6200 0.6750 0.8600 ;
        RECT  0.4050 1.7400 0.7150 1.8600 ;
        RECT  0.4050 0.7400 0.5250 1.8600 ;
        RECT  0.3600 0.8850 0.5250 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.7350 -0.1800 2.8550 0.7800 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.6150 1.7400 2.7350 2.7900 ;
        RECT  1.0150 2.2200 1.2550 2.7900 ;
        RECT  0.1650 1.5600 0.2850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.4150 1.7400 3.1550 1.7400 3.1550 1.8600 3.0350 1.8600 3.0350 1.6200 2.3350 1.6200
                 2.3350 2.2400 2.0550 2.2400 2.0550 2.1200 2.2150 2.1200 2.2150 1.5000 3.1550 1.5000
                 3.1550 1.6200 3.2950 1.6200 3.2950 0.7800 3.1550 0.7800 3.1550 0.5400 3.2750 0.5400
                 3.2750 0.6600 3.4150 0.6600 ;
        POLYGON  2.8550 1.0600 2.6150 1.0600 2.6150 1.0200 1.5750 1.0200 1.5750 1.5800 1.6750 1.5800
                 1.6750 1.8600 1.5550 1.8600 1.5550 1.7000 1.4550 1.7000 1.4550 0.6000 1.6950 0.6000
                 1.6950 0.7200 1.5750 0.7200 1.5750 0.9000 2.7350 0.9000 2.7350 0.9400 2.8550 0.9400 ;
        POLYGON  2.2150 0.7800 2.0950 0.7800 2.0950 0.4800 1.3350 0.4800 1.3350 1.1000 0.7650 1.1000
                 0.7650 1.5000 0.9550 1.5000 0.9550 1.5800 1.1400 1.5800 1.1400 1.9800 1.8150 1.9800
                 1.8150 1.8600 1.9750 1.8600 1.9750 1.7400 2.0950 1.7400 2.0950 1.9800 1.9350 1.9800
                 1.9350 2.1000 1.0200 2.1000 1.0200 1.7000 0.8350 1.7000 0.8350 1.6200 0.6450 1.6200
                 0.6450 0.9800 1.2150 0.9800 1.2150 0.3600 2.2150 0.3600 ;
    END
END XOR2X2

MACRO XOR2X1
    CLASS CORE ;
    FOREIGN XOR2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8550 1.2800 0.9750 1.5600 ;
        RECT  0.6800 1.4400 0.9750 1.5600 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 1.1800 2.8350 1.3000 ;
        RECT  2.0450 1.1800 2.3050 1.3800 ;
        RECT  1.9150 1.1400 2.1550 1.3000 ;
        RECT  1.3350 1.3600 1.5750 1.4800 ;
        RECT  1.4550 1.1800 1.5750 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 1.2950 0.2900 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.3950 -0.1800 2.5150 0.7800 ;
        RECT  0.4950 0.5500 0.7350 0.6700 ;
        RECT  0.6150 -0.1800 0.7350 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.2750 1.7400 2.3950 2.7900 ;
        RECT  0.5900 2.1600 0.8300 2.2800 ;
        RECT  0.5900 2.1600 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0750 1.7400 2.8150 1.7400 2.8150 1.8600 2.6950 1.8600 2.6950 1.6200 1.9550 1.6200
                 1.9550 2.2400 1.7150 2.2400 1.7150 2.1200 1.8350 2.1200 1.8350 1.5000 2.8150 1.5000
                 2.8150 1.6200 2.9550 1.6200 2.9550 0.7800 2.8150 0.7800 2.8150 0.5400 2.9350 0.5400
                 2.9350 0.6600 3.0750 0.6600 ;
        POLYGON  2.5150 1.0600 2.2750 1.0600 2.2750 1.0200 1.2150 1.0200 1.2150 1.6800 1.3100 1.6800
                 1.3100 1.8000 1.0700 1.8000 1.0700 1.6800 1.0950 1.6800 1.0950 0.6000 1.3350 0.6000
                 1.3350 0.7200 1.2150 0.7200 1.2150 0.9000 2.3950 0.9000 2.3950 0.9400 2.5150 0.9400 ;
        POLYGON  1.8750 0.7800 1.7550 0.7800 1.7550 0.4800 0.9750 0.4800 0.9750 1.1600 0.5500 1.1600
                 0.5500 1.2800 0.5300 1.2800 0.5300 1.9200 1.4750 1.9200 1.4750 1.8600 1.5500 1.8600
                 1.5500 1.7400 1.6700 1.7400 1.6700 1.9800 1.5950 1.9800 1.5950 2.0400 0.4100 2.0400
                 0.4100 1.0400 0.8550 1.0400 0.8550 0.3600 1.8750 0.3600 ;
    END
END XOR2X1

MACRO XNOR3XL
    CLASS CORE ;
    FOREIGN XNOR3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0800 1.3500 6.8100 1.4700 ;
        RECT  6.0800 1.2300 6.3650 1.4700 ;
        RECT  6.0800 0.9050 6.2000 1.4700 ;
        RECT  5.6950 0.9050 6.2000 1.0250 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2520  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.8450 0.9750 1.0250 1.3750 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.0700 0.3250 1.4700 ;
        RECT  0.0700 1.1750 0.3250 1.4350 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3704  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2700 1.5600 8.5100 2.2500 ;
        RECT  8.3900 0.3600 8.5100 2.2500 ;
        RECT  8.1350 0.6500 8.5100 0.8000 ;
        RECT  8.2700 0.3600 8.5100 0.8000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.7300 -0.1800 7.9700 0.3200 ;
        RECT  7.7900 -0.1800 7.9100 0.6700 ;
        RECT  1.8650 -0.1800 2.1050 0.3200 ;
        RECT  0.6850 -0.1800 0.9250 0.3200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.7300 2.2900 7.9700 2.7900 ;
        RECT  7.7900 1.6900 7.9100 2.7900 ;
        RECT  1.8650 2.2700 2.1050 2.7900 ;
        RECT  0.6850 2.2900 0.9250 2.7900 ;
        RECT  0.7450 1.9700 0.8650 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2300 1.3150 7.6700 1.3150 7.6700 2.1700 6.2600 2.1700 6.2600 1.8900 6.5600 1.8900
                 6.5600 2.0500 7.5500 2.0500 7.5500 0.6200 7.4200 0.6200 7.4200 0.4800 6.2600 0.4800
                 6.2600 0.3600 7.5400 0.3600 7.5400 0.5000 7.6700 0.5000 7.6700 1.1950 7.9900 1.1950
                 7.9900 1.0750 8.2300 1.0750 ;
        POLYGON  7.4300 0.8600 7.3450 0.8600 7.3450 1.8100 7.4300 1.8100 7.4300 1.9300 7.1900 1.9300
                 7.1900 1.8100 7.2250 1.8100 7.2250 0.8600 7.1900 0.8600 7.1900 0.7400 7.4300 0.7400 ;
        POLYGON  7.0500 1.7700 7.0400 1.7700 7.0400 1.7900 6.8000 1.7900 6.8000 1.7700 4.2750 1.7700
                 4.2750 1.6500 5.0950 1.6500 5.0950 0.7200 4.2700 0.7200 4.2700 0.6000 5.2150 0.6000
                 5.2150 1.6500 6.9300 1.6500 6.9300 0.7200 6.8000 0.7200 6.8000 0.6000 7.0500 0.6000 ;
        POLYGON  5.9600 0.7050 5.9000 0.7050 5.9000 0.7200 5.4800 0.7200 5.4800 1.4050 5.9600 1.4050
                 5.9600 1.5250 5.3600 1.5250 5.3600 0.6000 5.7200 0.6000 5.7200 0.5850 5.9600 0.5850 ;
        RECT  2.9850 1.8900 5.9600 2.0100 ;
        RECT  2.4050 0.3600 5.5550 0.4800 ;
        RECT  2.4050 2.1300 5.5550 2.2500 ;
        POLYGON  4.8400 1.0400 4.1700 1.0400 4.1700 1.4150 4.0500 1.4150 4.0500 0.9200 4.8400 0.9200 ;
        POLYGON  3.9850 0.7200 3.8400 0.7200 3.8400 1.7700 1.7250 1.7700 1.7250 2.1700 0.9850 2.1700
                 0.9850 1.8100 0.3250 1.8100 0.3250 1.9300 0.1450 1.9300 0.1450 1.6900 0.5050 1.6900
                 0.5050 0.9200 0.2050 0.9200 0.2050 0.4400 1.6050 0.4400 1.6050 0.3200 1.7250 0.3200
                 1.7250 0.5600 0.3250 0.5600 0.3250 0.8000 0.6250 0.8000 0.6250 1.6900 1.1050 1.6900
                 1.1050 2.0500 1.6050 2.0500 1.6050 1.6500 3.7200 1.6500 3.7200 0.6000 3.9850 0.6000 ;
        POLYGON  3.5850 1.0400 3.4050 1.0400 3.4050 1.0000 2.8100 1.0000 2.8100 1.1600 2.8850 1.1600
                 2.8850 1.2800 2.6450 1.2800 2.6450 1.1600 2.6900 1.1600 2.6900 0.8800 3.4050 0.8800
                 3.4050 0.8000 3.5850 0.8000 ;
        POLYGON  3.2250 1.5300 1.9400 1.5300 1.9400 0.6000 3.2050 0.6000 3.2050 0.7200 2.0600 0.7200
                 2.0600 1.4100 3.2250 1.4100 ;
        POLYGON  1.4850 1.4600 1.4050 1.4600 1.4050 1.8100 1.4650 1.8100 1.4650 1.9300 1.2250 1.9300
                 1.2250 1.8100 1.2850 1.8100 1.2850 1.4600 1.2450 1.4600 1.2450 1.3400 1.2850 1.3400
                 1.2850 0.8000 1.2250 0.8000 1.2250 0.6800 1.4650 0.6800 1.4650 0.8000 1.4050 0.8000
                 1.4050 1.3400 1.4850 1.3400 ;
    END
END XNOR3XL

MACRO XNOR3X1
    CLASS CORE ;
    FOREIGN XNOR3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4014  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2700 1.5600 8.5100 2.2500 ;
        RECT  8.3900 0.3600 8.5100 2.2500 ;
        RECT  8.1350 0.6500 8.5100 0.8000 ;
        RECT  8.2700 0.3600 8.5100 0.8000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0990  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.0700 0.3250 1.4700 ;
        RECT  0.0700 1.1750 0.3250 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2670  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.8400 1.0450 1.0250 1.3750 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0800 1.3500 6.8100 1.4700 ;
        RECT  6.0800 1.2300 6.3650 1.4700 ;
        RECT  6.0800 0.9050 6.2000 1.4700 ;
        RECT  5.7000 0.9050 6.2000 1.0250 ;
        END
    END C
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.7300 2.2900 7.9700 2.7900 ;
        RECT  7.7900 1.6900 7.9100 2.7900 ;
        RECT  1.8650 2.2700 2.1050 2.7900 ;
        RECT  0.6850 2.2900 0.9250 2.7900 ;
        RECT  0.7450 1.9700 0.8650 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.7300 -0.1800 7.9700 0.3200 ;
        RECT  7.7900 -0.1800 7.9100 0.6700 ;
        RECT  1.8650 -0.1800 2.1050 0.3200 ;
        RECT  0.6850 -0.1800 0.9250 0.3200 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  8.0700 1.3150 7.6700 1.3150 7.6700 2.1700 6.2600 2.1700 6.2600 1.8900 6.5600 1.8900
                 6.5600 2.0500 7.5500 2.0500 7.5500 0.6200 7.4200 0.6200 7.4200 0.4800 6.2600 0.4800
                 6.2600 0.3600 7.5400 0.3600 7.5400 0.5000 7.6700 0.5000 7.6700 1.1950 7.8300 1.1950
                 7.8300 1.0750 8.0700 1.0750 ;
        POLYGON  7.4300 0.8600 7.3450 0.8600 7.3450 1.8100 7.4300 1.8100 7.4300 1.9300 7.1900 1.9300
                 7.1900 1.8100 7.2250 1.8100 7.2250 0.8600 7.1900 0.8600 7.1900 0.7400 7.4300 0.7400 ;
        POLYGON  7.0500 1.7700 7.0400 1.7700 7.0400 1.7900 6.8000 1.7900 6.8000 1.7700 4.2750 1.7700
                 4.2750 1.6500 5.0950 1.6500 5.0950 0.7200 4.5250 0.7200 4.5250 0.6000 5.2150 0.6000
                 5.2150 1.6500 6.9300 1.6500 6.9300 0.7200 6.8000 0.7200 6.8000 0.6000 7.0500 0.6000 ;
        POLYGON  5.9600 0.7050 5.9000 0.7050 5.9000 0.7200 5.4800 0.7200 5.4800 1.4050 5.9600 1.4050
                 5.9600 1.5250 5.3600 1.5250 5.3600 0.6000 5.7200 0.6000 5.7200 0.5850 5.9600 0.5850 ;
        RECT  2.9850 1.8900 5.9600 2.0100 ;
        RECT  2.4050 0.3600 5.6400 0.4800 ;
        RECT  2.4050 2.1300 5.6400 2.2500 ;
        POLYGON  4.9700 1.0400 4.1700 1.0400 4.1700 1.2850 4.0500 1.2850 4.0500 0.9200 4.9700 0.9200 ;
        POLYGON  4.0750 0.7200 3.9300 0.7200 3.9300 1.7700 1.7250 1.7700 1.7250 2.1700 0.9850 2.1700
                 0.9850 1.8100 0.3250 1.8100 0.3250 1.9300 0.2050 1.9300 0.2050 1.6900 0.5050 1.6900
                 0.5050 0.9200 0.2050 0.9200 0.2050 0.4400 1.6050 0.4400 1.6050 0.3200 1.7250 0.3200
                 1.7250 0.5600 0.3250 0.5600 0.3250 0.8000 0.6250 0.8000 0.6250 1.6900 1.1050 1.6900
                 1.1050 2.0500 1.6050 2.0500 1.6050 1.6500 3.8100 1.6500 3.8100 0.6000 4.0750 0.6000 ;
        POLYGON  3.6900 1.0800 3.5700 1.0800 3.5700 1.0200 2.8100 1.0200 2.8100 1.1600 2.8850 1.1600
                 2.8850 1.2800 2.6450 1.2800 2.6450 1.1600 2.6900 1.1600 2.6900 0.9000 3.5700 0.9000
                 3.5700 0.8400 3.6900 0.8400 ;
        POLYGON  3.2250 1.5300 1.9400 1.5300 1.9400 0.6000 3.2050 0.6000 3.2050 0.7200 2.0600 0.7200
                 2.0600 1.4100 3.2250 1.4100 ;
        POLYGON  1.4850 1.5200 1.4050 1.5200 1.4050 1.8100 1.4650 1.8100 1.4650 1.9300 1.2250 1.9300
                 1.2250 1.8100 1.2850 1.8100 1.2850 1.5200 1.2450 1.5200 1.2450 1.4000 1.2850 1.4000
                 1.2850 0.8000 1.2250 0.8000 1.2250 0.6800 1.4650 0.6800 1.4650 0.8000 1.4050 0.8000
                 1.4050 1.4000 1.4850 1.4000 ;
    END
END XNOR3X1

MACRO XNOR2XL
    CLASS CORE ;
    FOREIGN XNOR2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7500 0.9800 0.8700 1.3400 ;
        RECT  0.6500 1.0800 0.8000 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9350 1.2400 2.8150 1.3600 ;
        RECT  2.0450 1.2300 2.3050 1.3800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1750 0.6200 0.2950 0.8850 ;
        RECT  0.1350 0.7650 0.2550 1.7600 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.4150 0.6800 2.6550 0.8000 ;
        RECT  2.4950 -0.1800 2.6150 0.8000 ;
        RECT  0.5950 -0.1800 0.7150 0.8600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3950 2.2200 2.6350 2.7900 ;
        RECT  0.6150 2.1600 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0550 2.0000 1.9950 2.0000 1.9950 2.1800 1.1750 2.1800 1.1750 2.0600 1.8750 2.0600
                 1.8750 1.8800 2.9350 1.8800 2.9350 1.1100 1.7950 1.1100 1.7950 1.2000 1.6750 1.2000
                 1.6750 0.9600 1.7950 0.9600 1.7950 0.9900 2.8950 0.9900 2.8950 0.6200 3.0150 0.6200
                 3.0150 0.8700 3.0550 0.8700 ;
        POLYGON  2.3750 0.4800 1.1950 0.4800 1.1950 0.6200 1.1350 0.6200 1.1350 1.5800 1.1550 1.5800
                 1.1550 1.7000 0.9150 1.7000 0.9150 1.5800 1.0150 1.5800 1.0150 0.5000 1.0750 0.5000
                 1.0750 0.3600 2.3750 0.3600 ;
        POLYGON  1.5550 1.9400 0.6750 1.9400 0.6750 1.6750 0.4100 1.6750 0.4100 1.2000 0.5300 1.2000
                 0.5300 1.5550 0.7950 1.5550 0.7950 1.8200 1.4350 1.8200 1.4350 0.6200 1.5550 0.6200 ;
    END
END XNOR2XL

MACRO XNOR2X4
    CLASS CORE ;
    FOREIGN XNOR2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.2100 2.2350 1.3450 ;
        RECT  1.7550 1.2100 2.0150 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7550 0.9000 3.8750 1.1400 ;
        RECT  3.2750 0.9700 3.8750 1.0900 ;
        RECT  3.4950 0.9400 3.8750 1.0900 ;
        RECT  2.5950 1.2100 3.3950 1.3300 ;
        RECT  3.2750 0.9700 3.3950 1.3300 ;
        RECT  3.0950 1.2100 3.3350 1.4100 ;
        RECT  2.5950 0.9300 2.7150 1.3300 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 1.7400 1.5750 2.2100 ;
        RECT  1.3950 0.6100 1.5150 0.8500 ;
        RECT  1.2750 1.7400 1.5750 1.8600 ;
        RECT  1.2750 1.3200 1.3950 1.8600 ;
        RECT  1.2150 0.7300 1.5150 0.8500 ;
        RECT  0.6500 0.8400 1.3350 0.9600 ;
        RECT  0.6500 1.3200 1.3950 1.4400 ;
        RECT  0.6500 1.1750 0.8000 1.4400 ;
        RECT  0.6500 0.7300 0.7700 1.5600 ;
        RECT  0.6150 1.4400 0.7350 2.2100 ;
        RECT  0.4950 0.7300 0.7700 0.8500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.4750 0.4200 3.7150 0.5400 ;
        RECT  3.4750 -0.1800 3.5950 0.5400 ;
        RECT  1.7550 0.5400 1.9950 0.6600 ;
        RECT  1.7550 -0.1800 1.8750 0.6600 ;
        RECT  0.9750 -0.1800 1.0950 0.7200 ;
        RECT  0.1350 -0.1800 0.2550 0.7200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.6550 1.7700 3.7750 2.7900 ;
        RECT  1.8150 2.0100 2.0550 2.1500 ;
        RECT  1.8150 2.0100 1.9350 2.7900 ;
        RECT  1.0350 1.5600 1.1550 2.7900 ;
        RECT  0.1950 1.5600 0.3150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.2550 1.9500 4.0150 1.9500 4.0150 0.7800 3.4200 0.7800 3.4200 0.8200 3.1550 0.8200
                 3.1550 1.0900 2.9150 1.0900 2.9150 0.9700 3.0350 0.9700 3.0350 0.7000 3.3000 0.7000
                 3.3000 0.6600 4.0150 0.6600 4.0150 0.5600 4.1350 0.5600 4.1350 1.8300 4.2550 1.8300 ;
        POLYGON  3.6350 1.6500 2.7750 1.6500 2.7750 2.0100 2.5350 2.0100 2.5350 1.6500 2.3550 1.6500
                 2.3550 0.6500 2.5950 0.6500 2.5950 0.7700 2.4750 0.7700 2.4750 1.5300 3.5150 1.5300
                 3.5150 1.2400 3.6350 1.2400 ;
        POLYGON  3.1350 2.2500 2.2200 2.2500 2.2200 1.8900 1.9550 1.8900 1.9550 1.6200 1.5150 1.6200
                 1.5150 1.2000 1.2550 1.2000 1.2550 1.0800 1.5150 1.0800 1.5150 0.9700 2.1150 0.9700
                 2.1150 0.4100 2.8950 0.4100 2.8950 0.4600 3.0150 0.4600 3.0150 0.5800 2.7750 0.5800
                 2.7750 0.5300 2.2350 0.5300 2.2350 1.0900 1.6350 1.0900 1.6350 1.5000 2.0750 1.5000
                 2.0750 1.7700 2.3400 1.7700 2.3400 2.1300 3.0150 2.1300 3.0150 1.7700 3.1350 1.7700 ;
    END
END XNOR2X4

MACRO XNOR2X2
    CLASS CORE ;
    FOREIGN XNOR2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.0600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.1100 1.7250 1.3800 ;
        RECT  1.4650 1.0200 1.7050 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.2600 3.5250 1.3800 ;
        RECT  2.6250 1.2300 2.8850 1.3800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8250 1.1750 1.0900 1.4350 ;
        RECT  0.6650 1.6200 0.9450 1.7400 ;
        RECT  0.8250 0.6800 0.9450 1.7400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.0600 0.1800 ;
        RECT  3.1250 0.7200 3.3650 0.8400 ;
        RECT  3.2050 -0.1800 3.3250 0.8400 ;
        RECT  1.2450 -0.1800 1.3650 0.7300 ;
        RECT  0.4050 -0.1800 0.5250 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.0600 2.7900 ;
        RECT  3.1250 1.7400 3.3650 1.8600 ;
        RECT  3.1250 1.7400 3.2450 2.7900 ;
        RECT  1.1450 2.1000 1.3850 2.2200 ;
        RECT  1.1450 2.1000 1.2650 2.7900 ;
        RECT  0.1850 2.1000 0.4250 2.2200 ;
        RECT  0.1850 2.1000 0.3050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.7650 1.6800 3.7250 1.6800 3.7250 1.8000 3.6050 1.8000 3.6050 1.6200 2.6550 1.6200
                 2.6550 2.2200 1.8850 2.2200 1.8850 2.1000 2.5350 2.1000 2.5350 1.5000 3.6450 1.5000
                 3.6450 1.1100 2.5050 1.1100 2.5050 1.2400 2.3850 1.2400 2.3850 0.9900 3.6050 0.9900
                 3.6050 0.6600 3.7250 0.6600 3.7250 0.8700 3.7650 0.8700 ;
        POLYGON  3.0850 0.5200 1.9050 0.5200 1.9050 0.6600 1.8450 0.6600 1.8450 0.7800 1.9650 0.7800
                 1.9650 1.7400 1.6250 1.7400 1.6250 1.6200 1.8450 1.6200 1.8450 0.9000 1.7250 0.9000
                 1.7250 0.5400 1.7850 0.5400 1.7850 0.4000 3.0850 0.4000 ;
        POLYGON  2.2650 1.9800 0.4250 1.9800 0.4250 1.3600 0.5450 1.3600 0.5450 1.2400 0.6650 1.2400
                 0.6650 1.4800 0.5450 1.4800 0.5450 1.8600 2.1450 1.8600 2.1450 0.6600 2.2650 0.6600 ;
    END
END XNOR2X2

MACRO XNOR2X1
    CLASS CORE ;
    FOREIGN XNOR2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.9350 1.3600 ;
        RECT  0.8150 1.1200 0.9350 1.3600 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6150 1.2600 2.8550 1.3800 ;
        RECT  1.9550 1.2800 2.7350 1.4000 ;
        RECT  2.0450 1.2300 2.3050 1.4000 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.8850 0.4550 1.0250 ;
        RECT  0.3350 0.6800 0.4550 1.0250 ;
        RECT  0.1350 0.8850 0.2550 2.1900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.4550 0.6800 2.6950 0.8000 ;
        RECT  2.5350 -0.1800 2.6550 0.8000 ;
        RECT  0.7550 -0.1800 0.8750 0.8600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3950 2.2400 2.6350 2.7900 ;
        RECT  0.6150 2.1800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0950 1.6600 3.0550 1.6600 3.0550 1.9000 1.9950 1.9000 1.9950 2.2000 1.1750 2.2000
                 1.1750 2.0800 1.8750 2.0800 1.8750 1.7800 2.9350 1.7800 2.9350 1.5400 2.9750 1.5400
                 2.9750 1.1100 1.7950 1.1100 1.7950 1.2200 1.6750 1.2200 1.6750 0.9800 1.7950 0.9800
                 1.7950 0.9900 2.9350 0.9900 2.9350 0.6200 3.0550 0.6200 3.0550 0.8700 3.0950 0.8700 ;
        POLYGON  2.4150 0.4800 1.2950 0.4800 1.2950 1.7200 0.9150 1.7200 0.9150 1.6000 1.1750 1.6000
                 1.1750 0.3600 2.4150 0.3600 ;
        POLYGON  1.7150 0.8600 1.5350 0.8600 1.5350 1.9600 0.6750 1.9600 0.6750 1.6750 0.4100 1.6750
                 0.4100 1.2200 0.5300 1.2200 0.5300 1.5550 0.7950 1.5550 0.7950 1.8400 1.4150 1.8400
                 1.4150 0.7400 1.5950 0.7400 1.5950 0.6200 1.7150 0.6200 ;
    END
END XNOR2X1

MACRO TLATXL
    CLASS CORE ;
    FOREIGN TLATXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0300 0.8500 1.4350 ;
        RECT  0.7300 1.0150 0.8500 1.4350 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.1400 3.4100 1.5900 ;
        RECT  3.2600 1.1400 3.3800 1.6150 ;
        END
    END G
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0100 0.5400 4.1300 0.7800 ;
        RECT  3.8400 1.4650 4.0800 1.7350 ;
        RECT  3.9600 0.6600 4.0800 1.7350 ;
        RECT  3.8100 1.6150 3.9300 1.8550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2400 0.6200 5.3600 1.1750 ;
        RECT  5.0400 1.0550 5.3600 1.1750 ;
        RECT  5.0400 1.0550 5.1600 1.7200 ;
        RECT  5.0000 1.1750 5.1600 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.8200 -0.1800 4.9400 0.8600 ;
        RECT  3.5900 -0.1800 3.7100 0.7800 ;
        RECT  2.3000 -0.1800 2.4200 0.3950 ;
        RECT  0.6150 -0.1800 0.7350 0.3950 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.6200 1.6000 4.7400 2.7900 ;
        RECT  3.3900 1.7350 3.5100 2.7900 ;
        RECT  1.9300 2.2150 2.1700 2.7900 ;
        RECT  0.5900 1.7950 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8800 1.3400 4.5000 1.3400 4.5000 1.6000 4.3200 1.6000 4.3200 1.7200 4.2000 1.7200
                 4.2000 1.4800 4.3800 1.4800 4.3800 1.1000 4.4000 1.1000 4.4000 0.6200 4.5200 0.6200
                 4.5200 1.2200 4.8800 1.2200 ;
        POLYGON  3.8400 1.0600 3.6000 1.0600 3.6000 1.0200 2.9000 1.0200 2.9000 1.5150 2.6500 1.5150
                 2.6500 1.8550 2.4100 1.8550 2.4100 1.7350 2.5300 1.7350 2.5300 1.5150 1.9300 1.5150
                 1.9300 1.3950 2.7800 1.3950 2.7800 0.6750 2.9000 0.6750 2.9000 0.9000 3.8400 0.9000 ;
        POLYGON  3.2900 0.7800 3.1700 0.7800 3.1700 0.5550 2.6600 0.5550 2.6600 0.6350 2.0100 0.6350
                 2.0100 0.6150 1.4300 0.6150 1.4300 1.4750 1.2100 1.4750 1.2100 1.5950 1.1100 1.5950
                 1.1100 2.0750 1.5200 2.0750 1.5200 1.9750 2.9700 1.9750 2.9700 1.7350 3.0900 1.7350
                 3.0900 2.0950 1.6400 2.0950 1.6400 2.1950 0.9900 2.1950 0.9900 1.6750 0.4100 1.6750
                 0.4100 1.3350 0.5300 1.3350 0.5300 1.5550 0.9900 1.5550 0.9900 1.3550 1.3100 1.3550
                 1.3100 0.4950 1.7100 0.4950 1.7100 0.3950 1.9500 0.3950 1.9500 0.4950 2.1300 0.4950
                 2.1300 0.5150 2.5400 0.5150 2.5400 0.4350 3.2900 0.4350 ;
        POLYGON  2.4900 1.2750 1.6700 1.2750 1.6700 1.8350 1.3500 1.8350 1.3500 1.9550 1.2300 1.9550
                 1.2300 1.7150 1.5500 1.7150 1.5500 0.7350 1.7900 0.7350 1.7900 0.8550 1.6700 0.8550
                 1.6700 1.1550 2.4900 1.1550 ;
        POLYGON  1.1900 1.2350 1.0700 1.2350 1.0700 0.8950 0.2900 0.8950 0.2900 1.9150 0.1700 1.9150
                 0.1700 0.9150 0.1350 0.9150 0.1350 0.6750 0.2550 0.6750 0.2550 0.7750 1.1900 0.7750 ;
    END
END TLATXL

MACRO TLATX4
    CLASS CORE ;
    FOREIGN TLATX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0450 0.5100 1.4400 ;
        RECT  0.3900 0.8350 0.5100 1.4400 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4800 1.4600 8.6300 1.7750 ;
        RECT  8.3250 1.4600 8.6300 1.7700 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1250 1.3200 2.2450 2.2100 ;
        RECT  1.2600 1.3200 2.2450 1.4400 ;
        RECT  1.0250 0.8000 2.1050 0.9200 ;
        RECT  1.9850 0.6800 2.1050 0.9200 ;
        RECT  1.2850 0.8000 1.4050 2.2100 ;
        RECT  1.2300 1.1750 1.4050 1.4350 ;
        RECT  1.0250 0.6800 1.1450 0.9200 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8250 0.8000 5.9450 0.9200 ;
        RECT  5.8250 0.6800 5.9450 0.9200 ;
        RECT  5.4850 1.3200 5.6050 2.2100 ;
        RECT  4.7100 1.3200 5.6050 1.4400 ;
        RECT  4.8650 0.6800 4.9850 0.9200 ;
        RECT  4.7100 1.1750 4.9450 1.5600 ;
        RECT  4.8250 0.8000 4.9450 1.5600 ;
        RECT  4.6450 1.4400 4.7650 2.2100 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        RECT  8.5450 -0.1800 8.6650 0.3800 ;
        RECT  7.2650 -0.1800 7.3850 0.4000 ;
        RECT  6.2450 -0.1800 6.4850 0.3200 ;
        RECT  5.2850 -0.1800 5.5250 0.3200 ;
        RECT  4.3250 -0.1800 4.5650 0.3200 ;
        RECT  3.3650 -0.1800 3.6050 0.3200 ;
        RECT  2.4050 -0.1800 2.6450 0.3200 ;
        RECT  1.4450 -0.1800 1.6850 0.3200 ;
        RECT  0.5450 -0.1800 0.6650 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        RECT  8.3850 1.9200 8.5050 2.7900 ;
        RECT  6.8050 1.8200 6.9250 2.7900 ;
        RECT  5.9050 1.5600 6.0250 2.7900 ;
        RECT  5.0650 1.5600 5.1850 2.7900 ;
        RECT  4.2250 1.5600 4.3450 2.7900 ;
        RECT  3.3850 1.5600 3.5050 2.7900 ;
        RECT  2.5450 1.5600 2.6650 2.7900 ;
        RECT  1.7050 1.5600 1.8250 2.7900 ;
        RECT  0.8650 1.5600 0.9850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.2050 0.8600 9.0850 0.8600 9.0850 1.3400 8.9250 1.3400 8.9250 2.0400 8.8050 2.0400
                 8.8050 1.3400 8.1250 1.3400 8.1250 1.5800 7.5850 1.5800 7.5850 1.7000 7.4650 1.7000
                 7.4650 1.4600 8.0050 1.4600 8.0050 1.2200 8.9650 1.2200 8.9650 0.7400 9.2050 0.7400 ;
        POLYGON  9.0450 0.5200 8.9250 0.5200 8.9250 0.6200 7.6450 0.6200 7.6450 0.6400 7.0250 0.6400
                 7.0250 0.5600 0.9050 0.5600 0.9050 0.6800 0.2550 0.6800 0.2550 0.9200 0.2400 0.9200
                 0.2400 1.5600 0.5050 1.5600 0.5050 1.8000 0.3850 1.8000 0.3850 1.6800 0.1200 1.6800
                 0.1200 0.8000 0.1350 0.8000 0.1350 0.5600 0.7850 0.5600 0.7850 0.4400 7.1450 0.4400
                 7.1450 0.5200 7.5250 0.5200 7.5250 0.5000 7.6450 0.5000 7.6450 0.4200 7.8850 0.4200
                 7.8850 0.5000 8.8050 0.5000 8.8050 0.4000 9.0450 0.4000 ;
        POLYGON  8.0250 0.8600 7.8850 0.8600 7.8850 1.3400 7.3450 1.3400 7.3450 1.8200 7.5850 1.8200
                 7.5850 1.8600 7.7050 1.8600 7.7050 1.9800 7.4650 1.9800 7.4650 1.9400 7.2250 1.9400
                 7.2250 1.7000 6.6250 1.7000 6.6250 1.3700 6.7450 1.3700 6.7450 1.5800 7.2250 1.5800
                 7.2250 1.2200 7.7650 1.2200 7.7650 0.7400 8.0250 0.7400 ;
        POLYGON  7.1050 1.4600 6.9850 1.4600 6.9850 1.2500 6.7850 1.2500 6.7850 1.2000 6.5050 1.2000
                 6.5050 2.2100 6.3850 2.2100 6.3850 1.2000 5.6250 1.2000 5.6250 1.0800 6.7850 1.0800
                 6.7850 0.6800 6.9050 0.6800 6.9050 1.1300 7.1050 1.1300 ;
        POLYGON  4.0250 0.9200 3.0650 0.9200 3.0650 1.0800 3.0850 1.0800 3.0850 1.3200 3.9250 1.3200
                 3.9250 2.2100 3.8050 2.2100 3.8050 1.4400 3.0850 1.4400 3.0850 2.2100 2.9650 2.2100
                 2.9650 1.2000 1.9250 1.2000 1.9250 1.0800 2.9450 1.0800 2.9450 0.6800 3.0650 0.6800
                 3.0650 0.8000 3.9050 0.8000 3.9050 0.6800 4.0250 0.6800 ;
    END
END TLATX4

MACRO TLATX2
    CLASS CORE ;
    FOREIGN TLATX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6200 0.6800 5.7400 2.1500 ;
        RECT  5.5800 1.1750 5.7400 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9400 0.8850 4.2800 1.1450 ;
        RECT  3.9400 0.6800 4.0600 2.1500 ;
        END
    END QN
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2050 1.4000 3.4650 1.6700 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.1250 0.8950 1.3550 ;
        RECT  0.5950 1.1250 0.8550 1.3800 ;
        END
    END D
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  6.0400 1.5000 6.1600 2.7900 ;
        RECT  5.2000 1.5000 5.3200 2.7900 ;
        RECT  4.3600 1.5000 4.4800 2.7900 ;
        RECT  3.5200 1.7900 3.6400 2.7900 ;
        RECT  2.0150 2.0800 2.2550 2.2000 ;
        RECT  2.0150 2.0800 2.1350 2.7900 ;
        RECT  0.6550 1.8200 0.7750 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  6.0400 -0.1800 6.1600 0.7300 ;
        RECT  5.2000 -0.1800 5.3200 0.7300 ;
        RECT  4.3600 -0.1800 4.4800 0.7300 ;
        RECT  3.4600 -0.1800 3.5800 0.4000 ;
        RECT  2.1750 -0.1800 2.2950 0.4000 ;
        RECT  0.5550 -0.1800 0.7950 0.3400 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  5.4600 1.3600 4.9000 1.3600 4.9000 2.1500 4.7800 2.1500 4.7800 0.6800 4.9000 0.6800
                 4.9000 1.2400 5.4600 1.2400 ;
        POLYGON  3.8200 1.2800 2.7750 1.2800 2.7750 1.5400 2.7350 1.5400 2.7350 1.7200 2.4950 1.7200
                 2.4950 1.5400 1.8150 1.5400 1.8150 1.4200 2.6550 1.4200 2.6550 0.6800 2.7750 0.6800
                 2.7750 1.1600 3.8200 1.1600 ;
        POLYGON  3.2800 1.9700 3.0400 1.9700 3.0400 1.9600 1.8950 1.9600 1.8950 2.1200 1.0150 2.1200
                 1.0150 1.6200 0.3550 1.6200 0.3550 1.3600 0.4750 1.3600 0.4750 1.5000 1.0150 1.5000
                 1.0150 1.3600 1.2950 1.3600 1.2950 0.5000 1.6950 0.5000 1.6950 0.4000 1.9350 0.4000
                 1.9350 0.5000 2.0150 0.5000 2.0150 0.5200 2.4150 0.5200 2.4150 0.4400 3.1650 0.4400
                 3.1650 0.9200 3.0450 0.9200 3.0450 0.5600 2.5350 0.5600 2.5350 0.6400 1.8950 0.6400
                 1.8950 0.6200 1.4150 0.6200 1.4150 1.6000 1.1350 1.6000 1.1350 2.0000 1.7750 2.0000
                 1.7750 1.8400 3.1600 1.8400 3.1600 1.8500 3.2800 1.8500 ;
        POLYGON  2.4950 1.3000 1.6550 1.3000 1.6550 1.8800 1.2550 1.8800 1.2550 1.7600 1.5350 1.7600
                 1.5350 0.7400 1.7750 0.7400 1.7750 0.8600 1.6550 0.8600 1.6550 1.1800 2.4950 1.1800 ;
        POLYGON  1.1750 1.2400 1.0550 1.2400 1.0550 1.0050 0.2350 1.0050 0.2350 1.7400 0.3550 1.7400
                 0.3550 1.9800 0.2350 1.9800 0.2350 1.8600 0.1150 1.8600 0.1150 0.8000 0.1350 0.8000
                 0.1350 0.6800 0.2550 0.6800 0.2550 0.8850 1.1750 0.8850 ;
    END
END TLATX2

MACRO TLATX1
    CLASS CORE ;
    FOREIGN TLATX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1150 0.8700 1.4350 ;
        RECT  0.6500 1.1100 0.8400 1.4350 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.0000 3.4100 1.4700 ;
        RECT  3.2600 1.0000 3.3800 1.5000 ;
        END
    END G
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9400 0.5900 4.0600 2.2100 ;
        RECT  3.8400 0.8850 4.0600 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.1700 0.6800 5.2900 2.1200 ;
        RECT  4.9450 0.9400 5.2900 1.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.7500 -0.1800 4.8700 0.7300 ;
        RECT  3.5200 -0.1800 3.6400 0.6400 ;
        RECT  2.2300 -0.1800 2.3500 0.3950 ;
        RECT  0.6150 -0.1800 0.7350 0.3950 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.7500 1.4700 4.8700 2.7900 ;
        RECT  3.5200 1.6200 3.6400 2.7900 ;
        RECT  1.9300 2.2150 2.1700 2.7900 ;
        RECT  0.5900 1.7950 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.0500 1.3300 4.4500 1.3300 4.4500 2.1200 4.3300 2.1200 4.3300 0.6800 4.4500 0.6800
                 4.4500 1.2100 5.0500 1.2100 ;
        POLYGON  3.7200 1.2200 3.6000 1.2200 3.6000 0.8800 2.8300 0.8800 2.8300 1.5150 2.6500 1.5150
                 2.6500 1.8550 2.4100 1.8550 2.4100 1.7350 2.5300 1.7350 2.5300 1.5150 1.9300 1.5150
                 1.9300 1.3950 2.7100 1.3950 2.7100 0.6750 2.8300 0.6750 2.8300 0.7600 3.7200 0.7600 ;
        POLYGON  3.2200 0.6400 3.1000 0.6400 3.1000 0.5550 2.5900 0.5550 2.5900 0.6350 1.9400 0.6350
                 1.9400 0.6150 1.4300 0.6150 1.4300 1.4750 1.2100 1.4750 1.2100 1.5950 1.1100 1.5950
                 1.1100 2.0750 1.5200 2.0750 1.5200 1.9750 3.0400 1.9750 3.0400 1.6800 3.1600 1.6800
                 3.1600 2.0950 1.6400 2.0950 1.6400 2.1950 0.9900 2.1950 0.9900 1.6750 0.4100 1.6750
                 0.4100 1.3350 0.5300 1.3350 0.5300 1.5550 0.9900 1.5550 0.9900 1.3550 1.3100 1.3550
                 1.3100 0.4950 1.7100 0.4950 1.7100 0.3950 1.9500 0.3950 1.9500 0.4950 2.0600 0.4950
                 2.0600 0.5150 2.4700 0.5150 2.4700 0.4350 3.1000 0.4350 3.1000 0.4000 3.2200 0.4000 ;
        POLYGON  2.4900 1.2750 1.6700 1.2750 1.6700 1.8350 1.3500 1.8350 1.3500 1.9550 1.2300 1.9550
                 1.2300 1.7150 1.5500 1.7150 1.5500 0.7350 1.7900 0.7350 1.7900 0.8550 1.6700 0.8550
                 1.6700 1.1550 2.4900 1.1550 ;
        POLYGON  1.1900 1.2350 1.0700 1.2350 1.0700 0.9900 0.2900 0.9900 0.2900 1.9150 0.1700 1.9150
                 0.1700 0.9150 0.1350 0.9150 0.1350 0.6750 0.2550 0.6750 0.2550 0.7950 0.2900 0.7950
                 0.2900 0.8700 1.1900 0.8700 ;
    END
END TLATX1

MACRO TLATSRXL
    CLASS CORE ;
    FOREIGN TLATSRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8850 1.2550 2.3050 1.4750 ;
        RECT  2.0450 1.2300 2.3050 1.4750 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7650 1.2700 2.8850 1.5950 ;
        RECT  2.6800 1.4550 2.8300 1.7250 ;
        END
    END G
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.1500 4.0450 1.4100 ;
        RECT  3.7650 1.1500 4.0450 1.3900 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5800 1.4650 5.9150 1.6100 ;
        RECT  5.7950 1.2600 5.9150 1.6100 ;
        RECT  5.5800 1.4650 5.7300 1.8150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 1.8300 ;
        RECT  1.2300 1.4650 1.4850 1.7250 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  5.9550 -0.1800 6.0750 0.7800 ;
        RECT  3.9850 0.4300 4.2250 0.5500 ;
        RECT  4.1050 -0.1800 4.2250 0.5500 ;
        RECT  1.7250 0.7400 1.9650 0.8600 ;
        RECT  1.7250 -0.1800 1.8450 0.8600 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  5.8750 2.2000 6.1150 2.7900 ;
        RECT  4.3650 2.0100 4.4850 2.7900 ;
        RECT  3.5250 2.2300 3.6450 2.7900 ;
        RECT  2.6850 2.2300 2.8050 2.7900 ;
        RECT  1.8450 2.2300 1.9650 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.5350 1.8400 6.4150 1.8400 6.4150 1.7200 6.3750 1.7200 6.3750 1.1400 5.5950 1.1400
                 5.5950 1.2000 5.4750 1.2000 5.4750 0.9600 5.5950 0.9600 5.5950 1.0200 6.3750 1.0200
                 6.3750 0.5400 6.4950 0.5400 6.4950 1.6000 6.5350 1.6000 ;
        POLYGON  6.4750 2.2200 6.2350 2.2200 6.2350 2.0800 5.5550 2.0800 5.5550 2.2200 5.3150 2.2200
                 5.3150 2.0800 4.9950 2.0800 4.9950 1.0400 4.8750 1.0400 4.8750 1.0300 3.4650 1.0300
                 3.4650 1.7100 3.1650 1.7100 3.1650 1.8300 3.0450 1.8300 3.0450 1.5900 3.3450 1.5900
                 3.3450 0.7200 3.2850 0.7200 3.2850 0.6000 3.5250 0.6000 3.5250 0.7200 3.4650 0.7200
                 3.4650 0.9100 5.1150 0.9100 5.1150 1.9600 6.3550 1.9600 6.3550 2.1000 6.4750 2.1000 ;
        POLYGON  5.3550 1.8400 5.2350 1.8400 5.2350 0.7900 3.6700 0.7900 3.6700 0.4800 2.9950 0.4800
                 2.9950 0.5400 2.2250 0.5400 2.2250 0.4200 2.8750 0.4200 2.8750 0.3600 3.7900 0.3600
                 3.7900 0.6700 5.2150 0.6700 5.2150 0.5400 5.3350 0.5400 5.3350 0.6600 5.3550 0.6600 ;
        POLYGON  4.8750 1.8000 4.7550 1.8000 4.7550 1.8900 3.8250 1.8900 3.8250 1.7700 4.6350 1.7700
                 4.6350 1.6800 4.8750 1.6800 ;
        POLYGON  4.2850 1.6500 3.7050 1.6500 3.7050 2.0700 2.7350 2.0700 2.7350 1.9650 2.2050 1.9650
                 2.2050 1.6050 2.4250 1.6050 2.4250 1.1100 1.7450 1.1100 1.7450 1.2600 1.6250 1.2600
                 1.6250 0.9900 2.4250 0.9900 2.4250 0.6800 2.5450 0.6800 2.5450 1.7250 2.3250 1.7250
                 2.3250 1.8450 2.8550 1.8450 2.8550 1.9500 3.5850 1.9500 3.5850 1.5300 4.1650 1.5300
                 4.1650 1.2700 4.2850 1.2700 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END TLATSRXL

MACRO TLATSRX4
    CLASS CORE ;
    FOREIGN TLATSRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7084  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.4900 2.5750 1.6100 ;
        RECT  2.3350 1.3150 2.5350 1.6100 ;
        RECT  2.4150 0.6200 2.5350 1.6100 ;
        RECT  1.4950 1.3150 2.5350 1.4350 ;
        RECT  1.4550 1.1750 1.6700 1.3150 ;
        RECT  1.3750 1.4900 1.6150 1.6100 ;
        RECT  1.4950 1.1750 1.6150 1.6100 ;
        RECT  1.4550 0.6200 1.5750 1.3150 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.8000 1.0750 10.9500 1.4350 ;
        RECT  10.7650 1.0300 10.8850 1.3900 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.1550 0.5650 1.3800 ;
        RECT  0.3250 1.1000 0.5650 1.3800 ;
        END
    END G
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7750 0.3600 9.0150 0.4800 ;
        RECT  8.1750 0.6900 8.8950 0.8100 ;
        RECT  8.7750 0.3600 8.8950 0.8100 ;
        RECT  8.1750 0.3800 8.2950 0.8100 ;
        RECT  7.2150 0.3800 8.2950 0.5000 ;
        RECT  6.6150 0.6900 7.3350 0.8100 ;
        RECT  7.2150 0.3800 7.3350 0.8100 ;
        RECT  6.6150 0.3800 6.7350 0.8100 ;
        RECT  6.1350 0.3800 6.7350 0.5000 ;
        RECT  5.5350 0.6900 6.2550 0.8100 ;
        RECT  6.1350 0.3800 6.2550 0.8100 ;
        RECT  5.5350 0.3800 5.6550 0.8100 ;
        RECT  5.0550 0.3800 5.6550 0.5000 ;
        RECT  4.5750 0.7900 5.1750 0.9100 ;
        RECT  5.0550 0.3800 5.1750 0.9100 ;
        RECT  4.5750 0.3800 4.6950 0.9100 ;
        RECT  4.0950 0.3800 4.6950 0.5000 ;
        RECT  3.6150 0.7900 4.2150 0.9100 ;
        RECT  4.0950 0.3800 4.2150 0.9100 ;
        RECT  3.6150 0.3800 3.7350 0.9100 ;
        RECT  3.1350 0.3800 3.7350 0.5000 ;
        RECT  2.6550 0.7900 3.2550 0.9100 ;
        RECT  3.1350 0.3800 3.2550 0.9100 ;
        RECT  2.6550 0.3800 2.7750 0.9100 ;
        RECT  2.1750 0.3800 2.7750 0.5000 ;
        RECT  1.6950 0.7900 2.2950 0.9100 ;
        RECT  2.1750 0.3800 2.2950 0.9100 ;
        RECT  1.6950 0.3800 1.8150 0.9100 ;
        RECT  1.2150 0.3800 1.8150 0.5000 ;
        RECT  0.9250 0.9600 1.3350 1.0800 ;
        RECT  1.2150 0.3800 1.3350 1.0800 ;
        RECT  0.9400 0.8850 1.0900 1.1450 ;
        RECT  0.9250 0.9600 1.0450 1.2000 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2150 1.1700 8.4550 1.2900 ;
        RECT  7.2650 1.2400 8.3350 1.3600 ;
        RECT  7.2650 1.1700 7.5250 1.3800 ;
        RECT  7.0550 1.1700 7.5250 1.2900 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7256  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.2150 0.9300 6.4950 1.0500 ;
        RECT  6.3750 0.6200 6.4950 1.0500 ;
        RECT  6.1750 1.4900 6.4150 1.6100 ;
        RECT  6.1750 1.3150 6.3350 1.6100 ;
        RECT  6.2150 0.9300 6.3350 1.6100 ;
        RECT  5.2900 1.3150 6.3350 1.4350 ;
        RECT  5.2150 1.4900 5.4550 1.6100 ;
        RECT  5.2900 1.3150 5.4550 1.6100 ;
        RECT  5.2900 1.1750 5.4400 1.6100 ;
        RECT  5.2950 0.6200 5.4150 1.6100 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  10.7050 0.5500 10.9450 0.6700 ;
        RECT  10.7050 -0.1800 10.8250 0.6700 ;
        RECT  8.4150 0.4500 8.6550 0.5700 ;
        RECT  8.5350 -0.1800 8.6550 0.5700 ;
        RECT  6.8550 0.4500 7.0950 0.5700 ;
        RECT  6.9750 -0.1800 7.0950 0.5700 ;
        RECT  5.7750 0.4500 6.0150 0.5700 ;
        RECT  5.8950 -0.1800 6.0150 0.5700 ;
        RECT  4.8150 -0.1800 4.9350 0.6700 ;
        RECT  3.8550 -0.1800 3.9750 0.6700 ;
        RECT  2.8950 -0.1800 3.0150 0.6700 ;
        RECT  1.9350 -0.1800 2.0550 0.6700 ;
        RECT  0.9750 -0.1800 1.0950 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  10.9250 1.7950 11.0450 2.7900 ;
        RECT  9.2950 2.2300 9.5350 2.7900 ;
        RECT  8.5150 2.2300 8.6350 2.7900 ;
        RECT  7.6750 2.2300 7.7950 2.7900 ;
        RECT  6.6550 1.9800 6.8950 2.1000 ;
        RECT  6.6550 1.9800 6.7750 2.7900 ;
        RECT  5.6950 1.9700 5.9350 2.0900 ;
        RECT  5.6950 1.9700 5.8150 2.7900 ;
        RECT  4.7350 1.9700 4.9750 2.0900 ;
        RECT  4.7350 1.9700 4.8550 2.7900 ;
        RECT  3.7750 1.9700 4.0150 2.0900 ;
        RECT  3.7750 1.9700 3.8950 2.7900 ;
        RECT  2.8150 1.9700 3.0550 2.0900 ;
        RECT  2.8150 1.9700 2.9350 2.7900 ;
        RECT  1.8550 1.9700 2.0950 2.0900 ;
        RECT  1.8550 1.9700 1.9750 2.7900 ;
        RECT  0.9550 2.0700 1.0750 2.7900 ;
        RECT  0.1350 1.5500 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.4650 1.9150 11.3450 1.9150 11.3450 0.9100 10.3100 0.9100 10.3100 0.8100
                 10.0450 0.8100 10.0450 0.4800 9.9250 0.4800 9.9250 0.3600 10.1650 0.3600
                 10.1650 0.6900 10.4300 0.6900 10.4300 0.7900 11.2450 0.7900 11.2450 0.6200
                 11.3650 0.6200 11.3650 0.7400 11.4650 0.7400 ;
        POLYGON  11.2050 1.6750 10.6450 1.6750 10.6450 2.1550 10.0450 2.1550 10.0450 2.1100
                 7.7100 2.1100 7.7100 1.8600 6.3850 1.8600 6.3850 1.8500 0.5550 1.8500 0.5550 1.5000
                 0.6850 1.5000 0.6850 0.9800 0.2750 0.9800 0.2750 0.6200 0.3950 0.6200 0.3950 0.8600
                 0.8050 0.8600 0.8050 1.7300 6.5050 1.7300 6.5050 1.7400 7.8300 1.7400 7.8300 1.9900
                 10.0450 1.9900 10.0450 1.6300 9.5450 1.6300 9.5450 1.1700 9.6650 1.1700 9.6650 1.5100
                 10.1650 1.5100 10.1650 2.0350 10.5250 2.0350 10.5250 1.1500 10.1450 1.1500
                 10.1450 1.0300 10.6450 1.0300 10.6450 1.5550 11.0850 1.5550 11.0850 1.3350
                 11.2050 1.3350 ;
        POLYGON  10.4050 1.9150 10.2850 1.9150 10.2850 1.3900 9.9050 1.3900 9.9050 1.0500 8.0950 1.0500
                 8.0950 1.1200 7.8550 1.1200 7.8550 0.9300 9.7050 0.9300 9.7050 0.6200 9.8250 0.6200
                 9.8250 0.9300 10.0250 0.9300 10.0250 1.2700 10.4050 1.2700 ;
        RECT  8.8150 1.7500 9.9250 1.8700 ;
        POLYGON  9.2150 1.4300 8.6950 1.4300 8.6950 1.6200 8.1550 1.6200 8.1550 1.8700 8.0350 1.8700
                 8.0350 1.6200 6.8150 1.6200 6.8150 1.2900 6.4550 1.2900 6.4550 1.1700 6.8150 1.1700
                 6.8150 0.9300 7.6150 0.9300 7.6150 0.6200 7.7350 0.6200 7.7350 1.0500 6.9350 1.0500
                 6.9350 1.5000 8.0350 1.5000 8.0350 1.4800 8.1550 1.4800 8.1550 1.5000 8.5750 1.5000
                 8.5750 1.3100 9.2150 1.3100 ;
        POLYGON  4.4950 1.6100 4.2550 1.6100 4.2550 1.4900 4.3350 1.4900 4.3350 1.1500 3.4950 1.1500
                 3.4950 1.4900 3.5350 1.4900 3.5350 1.6100 3.2950 1.6100 3.2950 1.4900 3.3750 1.4900
                 3.3750 1.1500 2.6550 1.1500 2.6550 1.0300 3.3750 1.0300 3.3750 0.6200 3.4950 0.6200
                 3.4950 1.0300 4.3350 1.0300 4.3350 0.6200 4.4550 0.6200 4.4550 1.4900 4.4950 1.4900 ;
    END
END TLATSRX4

MACRO TLATSRX2
    CLASS CORE ;
    FOREIGN TLATSRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 1.0100 3.7000 1.4800 ;
        RECT  3.5650 0.9800 3.6850 1.4800 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.1600 0.8350 1.5800 ;
        RECT  0.6500 1.1600 0.8350 1.5650 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.3300 3.1200 1.7250 ;
        RECT  2.8800 1.3300 3.1200 1.4500 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6250 1.2150 4.9150 1.4300 ;
        RECT  4.6250 1.0950 4.7450 1.4700 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5250 0.9400 5.7850 1.0900 ;
        RECT  5.2850 0.9400 5.7850 1.0600 ;
        RECT  5.2850 0.6150 5.4050 1.3350 ;
        RECT  5.1850 1.2150 5.3050 2.1100 ;
        RECT  5.1850 0.4950 5.3050 0.7350 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8850 0.8850 7.1800 1.1450 ;
        RECT  6.8850 0.7650 7.0050 1.5800 ;
        RECT  6.8650 1.4600 6.9850 2.1100 ;
        RECT  6.8650 0.5950 6.9850 0.8850 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  7.2850 -0.1800 7.4050 0.6450 ;
        RECT  6.4450 -0.1800 6.5650 0.6450 ;
        RECT  5.6050 -0.1800 5.7250 0.6450 ;
        RECT  4.7650 -0.1800 4.8850 0.7350 ;
        RECT  2.7150 0.6100 2.9550 0.7300 ;
        RECT  2.8350 -0.1800 2.9550 0.7300 ;
        RECT  0.4950 0.6800 0.7350 0.8000 ;
        RECT  0.4950 -0.1800 0.6150 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  7.2850 1.4600 7.4050 2.7900 ;
        RECT  6.4450 1.4600 6.5650 2.7900 ;
        RECT  5.6050 1.4600 5.7250 2.7900 ;
        RECT  4.7650 1.5900 4.8850 2.7900 ;
        RECT  3.8650 2.2300 3.9850 2.7900 ;
        RECT  3.1450 2.2300 3.2650 2.7900 ;
        RECT  2.2450 2.2900 2.4850 2.7900 ;
        RECT  0.7150 1.9400 0.8350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.7650 1.2400 6.1450 1.2400 6.1450 2.1100 6.0250 2.1100 6.0250 0.5950 6.1450 0.5950
                 6.1450 1.1200 6.7650 1.1200 ;
        POLYGON  5.1650 1.0950 4.9250 1.0950 4.9250 0.9750 4.4650 0.9750 4.4650 2.1100 4.3450 2.1100
                 4.3450 0.9750 4.1250 0.9750 4.1250 0.5000 3.1950 0.5000 3.1950 0.9700 2.2750 0.9700
                 2.2750 0.4800 2.1550 0.4800 2.1550 0.3600 2.3950 0.3600 2.3950 0.8500 3.0750 0.8500
                 3.0750 0.3800 4.2450 0.3800 4.2450 0.8550 5.1650 0.8550 ;
        POLYGON  4.1850 2.1100 2.4100 2.1100 2.4100 2.1700 1.4950 2.1700 1.4950 1.7500 1.6150 1.7500
                 1.6150 1.5700 1.6550 1.5700 1.6550 0.6200 1.7750 0.6200 1.7750 1.6900 1.7350 1.6900
                 1.7350 1.8700 1.6150 1.8700 1.6150 2.0500 2.2900 2.0500 2.2900 1.9900 4.0650 1.9900
                 4.0650 1.2700 4.1850 1.2700 ;
        POLYGON  3.9400 1.7200 3.6250 1.7200 3.6250 1.8400 3.5050 1.8400 3.5050 1.7200 3.2400 1.7200
                 3.2400 1.2100 1.9150 1.2100 1.9150 0.5000 1.5350 0.5000 1.5350 1.4500 1.4150 1.4500
                 1.4150 1.0400 0.5150 1.0400 0.5150 1.2000 0.3950 1.2000 0.3950 0.9200 1.4150 0.9200
                 1.4150 0.3800 2.0350 0.3800 2.0350 0.9600 2.0950 0.9600 2.0950 1.0900 3.3600 1.0900
                 3.3600 1.6000 3.8200 1.6000 3.8200 0.8600 3.4750 0.8600 3.4750 0.6200 3.5950 0.6200
                 3.5950 0.7400 3.9400 0.7400 ;
        POLYGON  2.8450 1.8700 2.0950 1.8700 2.0950 1.9300 1.8550 1.9300 1.8550 1.8100 1.9750 1.8100
                 1.9750 1.7500 2.8450 1.7500 ;
        POLYGON  1.2350 1.2800 1.0750 1.2800 1.0750 1.8200 0.3550 1.8200 0.3550 1.9900 0.2350 1.9900
                 0.2350 1.8700 0.1550 1.8700 0.1550 0.8600 0.1350 0.8600 0.1350 0.6200 0.2550 0.6200
                 0.2550 0.7400 0.2750 0.7400 0.2750 1.7000 0.9550 1.7000 0.9550 1.1600 1.2350 1.1600 ;
    END
END TLATSRX2

MACRO TLATSRX1
    CLASS CORE ;
    FOREIGN TLATSRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.5200 ;
        RECT  1.9450 1.2600 2.2500 1.4300 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.2000 3.0050 1.4500 ;
        RECT  2.6250 1.2000 2.8850 1.4700 ;
        END
    END G
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4950 1.1600 3.8450 1.4100 ;
        RECT  3.4950 1.1400 3.7550 1.4100 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5800 1.2800 5.8350 1.7350 ;
        RECT  5.7150 1.2600 5.8350 1.7350 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2888  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 0.9200 ;
        RECT  1.2850 0.8000 1.4050 2.2100 ;
        RECT  1.2300 1.4650 1.4050 1.7250 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  5.9550 -0.1800 6.0750 0.7800 ;
        RECT  4.0250 0.4200 4.2650 0.5400 ;
        RECT  4.1450 -0.1800 4.2650 0.5400 ;
        RECT  1.7850 -0.1800 1.9050 0.7300 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  5.8750 2.2000 6.1150 2.7900 ;
        RECT  4.3050 2.0100 4.4250 2.7900 ;
        RECT  3.4650 2.2300 3.5850 2.7900 ;
        RECT  2.6050 2.2300 2.7250 2.7900 ;
        RECT  1.7050 1.5900 1.8250 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.5350 1.8400 6.4150 1.8400 6.4150 1.7200 6.3750 1.7200 6.3750 1.0200 5.5950 1.0200
                 5.5950 1.1400 5.4750 1.1400 5.4750 0.9000 6.3750 0.9000 6.3750 0.5400 6.4950 0.5400
                 6.4950 1.6000 6.5350 1.6000 ;
        POLYGON  6.4750 2.2200 6.2350 2.2200 6.2350 2.0800 5.5550 2.0800 5.5550 2.2200 5.3150 2.2200
                 5.3150 2.0800 4.9950 2.0800 4.9950 1.0400 4.8750 1.0400 4.8750 1.0200 3.3750 1.0200
                 3.3750 1.7100 3.1050 1.7100 3.1050 1.8300 2.9850 1.8300 2.9850 1.5900 3.2550 1.5900
                 3.2550 0.6000 3.5650 0.6000 3.5650 0.7200 3.3750 0.7200 3.3750 0.9000 5.1150 0.9000
                 5.1150 1.9600 6.3550 1.9600 6.3550 2.1000 6.4750 2.1000 ;
        POLYGON  5.3550 1.8400 5.2350 1.8400 5.2350 0.7800 3.7300 0.7800 3.7300 0.4800 2.7900 0.4800
                 2.7900 0.5400 2.2850 0.5400 2.2850 0.4200 2.6700 0.4200 2.6700 0.3600 3.8500 0.3600
                 3.8500 0.6600 5.2150 0.6600 5.2150 0.5400 5.3350 0.5400 5.3350 0.6600 5.3550 0.6600 ;
        POLYGON  4.8750 1.8000 4.7550 1.8000 4.7550 1.8900 3.7650 1.8900 3.7650 1.7700 4.6350 1.7700
                 4.6350 1.6800 4.8750 1.6800 ;
        POLYGON  4.2250 1.6500 3.6450 1.6500 3.6450 2.0700 2.1250 2.0700 2.1250 1.6400 2.3700 1.6400
                 2.3700 1.0550 1.7250 1.0550 1.7250 1.2600 1.6050 1.2600 1.6050 0.9350 2.4850 0.9350
                 2.4850 0.6800 2.6050 0.6800 2.6050 1.0550 2.4900 1.0550 2.4900 1.7600 2.2450 1.7600
                 2.2450 1.9500 3.5250 1.9500 3.5250 1.5300 4.1050 1.5300 4.1050 1.2700 4.2250 1.2700 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END TLATSRX1

MACRO TLATNXL
    CLASS CORE ;
    FOREIGN TLATNXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7200 1.0400 0.8400 1.4200 ;
        RECT  0.6500 1.0650 0.8000 1.4350 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.2750 3.4100 1.7250 ;
        RECT  3.2900 1.2500 3.4100 1.7250 ;
        END
    END GN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9300 1.5850 4.0500 2.0900 ;
        RECT  3.8400 1.3450 3.9900 1.7250 ;
        RECT  3.8100 0.6400 3.9300 1.4650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.1600 1.4350 5.2800 1.6750 ;
        RECT  5.0000 1.1750 5.1600 1.4350 ;
        RECT  5.0400 0.5750 5.1600 1.5550 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.6200 -0.1800 4.7400 0.8150 ;
        RECT  3.3300 -0.1800 3.4500 0.8800 ;
        RECT  2.0400 -0.1800 2.1600 0.6400 ;
        RECT  0.6500 -0.1800 0.7700 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.7400 1.5550 4.8600 2.7900 ;
        RECT  3.5100 1.9700 3.6300 2.7900 ;
        RECT  2.3000 2.0800 2.4200 2.7900 ;
        RECT  0.6150 2.0800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8800 1.0750 4.4400 1.0750 4.4400 1.6750 4.3200 1.6750 4.3200 0.9550 4.2000 0.9550
                 4.2000 0.5750 4.3200 0.5750 4.3200 0.8350 4.4400 0.8350 4.4400 0.9550 4.8800 0.9550 ;
        POLYGON  3.8100 0.4800 3.6900 0.4800 3.6900 1.1200 3.0900 1.1200 3.0900 0.5200 2.7300 0.5200
                 2.7300 1.4800 2.9000 1.4800 2.9000 1.7200 2.7800 1.7200 2.7800 1.6000 2.6100 1.6000
                 2.6100 1.2400 2.2700 1.2400 2.2700 1.3600 2.1500 1.3600 2.1500 1.1200 2.6100 1.1200
                 2.6100 0.6400 2.4600 0.6400 2.4600 0.4000 3.2100 0.4000 3.2100 1.0000 3.5700 1.0000
                 3.5700 0.3600 3.8100 0.3600 ;
        POLYGON  3.2100 2.1100 3.0900 2.1100 3.0900 1.9900 3.0200 1.9900 3.0200 1.9650 2.5600 1.9650
                 2.5600 1.9600 1.3600 1.9600 1.3600 0.9200 0.5300 0.9200 0.5300 0.9800 0.4100 0.9800
                 0.4100 0.7400 0.5300 0.7400 0.5300 0.8000 1.4800 0.8000 1.4800 1.2200 1.6700 1.2200
                 1.6700 1.1000 1.7900 1.1000 1.7900 1.3400 1.4800 1.3400 1.4800 1.8400 2.6800 1.8400
                 2.6800 1.8450 3.0200 1.8450 3.0200 1.3600 2.8500 1.3600 2.8500 0.6400 2.9700 0.6400
                 2.9700 1.2400 3.1400 1.2400 3.1400 1.8450 3.2100 1.8450 ;
        POLYGON  2.4900 1.0000 2.3700 1.0000 2.3700 0.9800 2.0300 0.9800 2.0300 1.5800 1.7200 1.5800
                 1.7200 1.7000 1.6000 1.7000 1.6000 1.4600 1.9100 1.4600 1.9100 0.9800 1.6000 0.9800
                 1.6000 0.6800 1.2900 0.6800 1.2900 0.4000 1.4100 0.4000 1.4100 0.5600 1.7200 0.5600
                 1.7200 0.8600 2.3700 0.8600 2.3700 0.7600 2.4900 0.7600 ;
        POLYGON  1.2400 1.3000 1.1200 1.3000 1.1200 1.6750 0.2550 1.6750 0.2550 1.7950 0.1350 1.7950
                 0.1350 1.5550 0.1700 1.5550 0.1700 0.4000 0.2900 0.4000 0.2900 1.5550 1.0000 1.5550
                 1.0000 1.1800 1.2400 1.1800 ;
    END
END TLATNXL

MACRO TLATNX4
    CLASS CORE ;
    FOREIGN TLATNX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 0.9300 0.8550 1.1400 ;
        RECT  0.5550 1.0200 0.7950 1.2000 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7700 1.3450 8.9200 1.7600 ;
        RECT  8.7950 1.1200 8.9150 1.7600 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2950 1.3200 2.4150 2.2100 ;
        RECT  1.5200 1.3200 2.4150 1.4400 ;
        RECT  1.0950 0.8000 2.1750 0.9200 ;
        RECT  2.0550 0.6800 2.1750 0.9200 ;
        RECT  1.5500 0.8000 1.6700 1.5600 ;
        RECT  1.4550 1.4400 1.5750 2.2100 ;
        RECT  1.5200 1.1750 1.6700 1.5600 ;
        RECT  1.0950 0.6800 1.2150 0.9200 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9350 0.8000 6.0150 0.9200 ;
        RECT  5.8950 0.6800 6.0150 0.9200 ;
        RECT  5.6550 1.5200 5.7750 2.2100 ;
        RECT  4.9450 1.5200 5.7750 1.6400 ;
        RECT  4.8150 1.5500 5.2050 1.6700 ;
        RECT  5.0850 0.8000 5.2050 1.6700 ;
        RECT  4.9350 0.6800 5.0550 0.9200 ;
        RECT  4.8150 1.5500 4.9350 2.2100 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.7350 -0.1800 8.8550 0.4000 ;
        RECT  7.3350 -0.1800 7.4550 0.4000 ;
        RECT  6.3150 -0.1800 6.5550 0.3200 ;
        RECT  5.3550 -0.1800 5.5950 0.3200 ;
        RECT  4.3950 -0.1800 4.6350 0.3200 ;
        RECT  3.4350 -0.1800 3.6750 0.3200 ;
        RECT  2.4750 -0.1800 2.7150 0.3200 ;
        RECT  1.5150 -0.1800 1.7550 0.3200 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.7550 1.8800 8.8750 2.7900 ;
        RECT  6.9150 1.6600 7.1550 2.0600 ;
        RECT  6.9150 1.6600 7.0350 2.7900 ;
        RECT  6.0750 1.5600 6.1950 2.7900 ;
        RECT  5.2350 1.7900 5.3550 2.7900 ;
        RECT  4.3950 1.5600 4.5150 2.7900 ;
        RECT  3.5550 1.5600 3.6750 2.7900 ;
        RECT  2.7150 1.5600 2.8350 2.7900 ;
        RECT  1.8750 1.5600 1.9950 2.7900 ;
        RECT  1.0350 1.5600 1.1550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.4550 0.8600 9.3350 0.8600 9.3350 1.0000 9.2950 1.0000 9.2950 2.0000 9.1750 2.0000
                 9.1750 1.0000 8.6350 1.0000 8.6350 1.4000 8.3950 1.4000 8.3950 0.8800 9.2150 0.8800
                 9.2150 0.7400 9.4550 0.7400 ;
        POLYGON  9.2350 0.5200 9.0950 0.5200 9.0950 0.6400 8.4950 0.6400 8.4950 0.6200 7.8550 0.6200
                 7.8550 1.5000 7.9750 1.5000 7.9750 1.6200 7.7350 1.6200 7.7350 0.6400 7.0950 0.6400
                 7.0950 0.5600 0.9750 0.5600 0.9750 0.6800 0.2550 0.6800 0.2550 1.3200 0.5750 1.3200
                 0.5750 1.8000 0.4550 1.8000 0.4550 1.4400 0.1350 1.4400 0.1350 0.5600 0.8550 0.5600
                 0.8550 0.4400 7.2150 0.4400 7.2150 0.5200 7.7350 0.5200 7.7350 0.5000 8.1350 0.5000
                 8.1350 0.4000 8.3750 0.4000 8.3750 0.5000 8.6150 0.5000 8.6150 0.5200 8.9750 0.5200
                 8.9750 0.4000 9.2350 0.4000 ;
        POLYGON  8.2150 2.0000 8.0950 2.0000 8.0950 1.8600 7.4950 1.8600 7.4950 1.5000 6.8150 1.5000
                 6.8150 1.2600 6.9350 1.2600 6.9350 1.3800 7.6150 1.3800 7.6150 1.7400 8.0950 1.7400
                 8.0950 0.8600 7.9750 0.8600 7.9750 0.7400 8.2150 0.7400 ;
        POLYGON  7.5550 1.2600 7.4350 1.2600 7.4350 1.1400 6.6750 1.1400 6.6750 2.1200 6.5550 2.1200
                 6.5550 1.2600 5.6950 1.2600 5.6950 1.1400 6.5550 1.1400 6.5550 1.0200 6.8550 1.0200
                 6.8550 0.6800 6.9750 0.6800 6.9750 1.0200 7.5550 1.0200 ;
        POLYGON  4.0950 0.9200 3.2550 0.9200 3.2550 1.3200 4.0950 1.3200 4.0950 2.2100 3.9750 2.2100
                 3.9750 1.4400 3.2550 1.4400 3.2550 2.2100 3.1350 2.2100 3.1350 1.2000 2.0950 1.2000
                 2.0950 1.0800 3.1350 1.0800 3.1350 0.9200 3.0150 0.9200 3.0150 0.6800 3.1350 0.6800
                 3.1350 0.8000 3.9750 0.8000 3.9750 0.6800 4.0950 0.6800 ;
    END
END TLATNX4

MACRO TLATNX2
    CLASS CORE ;
    FOREIGN TLATNX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.4650 0.9400 5.7850 1.0900 ;
        RECT  5.4650 0.6400 5.5850 1.9900 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 0.8850 3.9900 1.1450 ;
        RECT  3.7850 0.6400 3.9050 1.9900 ;
        END
    END QN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 0.9400 3.1750 1.2100 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.0700 0.8750 1.1900 ;
        RECT  0.3050 1.2300 0.7150 1.3800 ;
        RECT  0.5950 1.0700 0.7150 1.3800 ;
        END
    END D
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.8850 1.3400 6.0050 2.7900 ;
        RECT  5.0450 1.3400 5.1650 2.7900 ;
        RECT  4.2050 1.3400 4.3250 2.7900 ;
        RECT  3.3050 1.4000 3.5450 1.6400 ;
        RECT  3.3050 1.4000 3.4250 2.7900 ;
        RECT  2.0550 2.2700 2.2950 2.7900 ;
        RECT  0.7350 1.8100 0.8550 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.8850 -0.1800 6.0050 0.6900 ;
        RECT  5.0450 -0.1800 5.1650 0.6900 ;
        RECT  4.2050 -0.1800 4.3250 0.6900 ;
        RECT  3.2450 -0.1800 3.4850 0.3400 ;
        RECT  2.0150 -0.1800 2.1350 0.7100 ;
        RECT  0.5550 -0.1800 0.6750 0.7100 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  5.3450 1.2000 4.7450 1.2000 4.7450 1.9900 4.6250 1.9900 4.6250 0.6400 4.7450 0.6400
                 4.7450 1.0800 5.3450 1.0800 ;
        POLYGON  3.6250 1.2000 3.5050 1.2000 3.5050 0.8200 3.2300 0.8200 3.2300 0.5800 2.5550 0.5800
                 2.5550 1.7900 2.7750 1.7900 2.7750 1.9100 2.4350 1.9100 2.4350 1.4300 2.1750 1.4300
                 2.1750 1.5500 2.0550 1.5500 2.0550 1.3100 2.4350 1.3100 2.4350 0.4600 3.3500 0.4600
                 3.3500 0.7000 3.6250 0.7000 ;
        POLYGON  3.0650 2.1500 1.1150 2.1500 1.1150 1.5500 1.5350 1.5500 1.5350 1.0700 1.0350 1.0700
                 1.0350 0.9500 0.4750 0.9500 0.4750 1.0700 0.3550 1.0700 0.3550 0.8300 1.6550 0.8300
                 1.6550 1.3500 1.6950 1.3500 1.6950 1.5900 1.6550 1.5900 1.6550 1.6700 1.2350 1.6700
                 1.2350 2.0300 2.9450 2.0300 2.9450 1.4600 2.6750 1.4600 2.6750 0.7000 3.0050 0.7000
                 3.0050 0.8200 2.7950 0.8200 2.7950 1.3400 3.0650 1.3400 ;
        POLYGON  2.3150 1.1500 1.9350 1.1500 1.9350 1.9100 1.3550 1.9100 1.3550 1.7900 1.8150 1.7900
                 1.8150 1.1500 1.7750 1.1500 1.7750 0.7100 1.1950 0.7100 1.1950 0.4700 1.3150 0.4700
                 1.3150 0.5900 1.8950 0.5900 1.8950 1.0300 2.3150 1.0300 ;
        POLYGON  1.4150 1.4300 0.9550 1.4300 0.9550 1.6200 0.4350 1.6200 0.4350 1.9300 0.3150 1.9300
                 0.3150 1.7400 0.0650 1.7400 0.0650 0.5900 0.1350 0.5900 0.1350 0.4700 0.2550 0.4700
                 0.2550 0.7100 0.1850 0.7100 0.1850 1.5000 0.8350 1.5000 0.8350 1.3100 1.4150 1.3100 ;
    END
END TLATNX2

MACRO TLATNX1
    CLASS CORE ;
    FOREIGN TLATNX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.4000 0.7600 1.5200 ;
        RECT  0.6400 1.0200 0.7600 1.5200 ;
        RECT  0.3600 1.0500 0.5100 1.5200 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1950 1.1650 3.4650 1.3800 ;
        RECT  3.1950 1.0900 3.3150 1.4700 ;
        END
    END GN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8400 1.1750 3.9900 1.4350 ;
        RECT  3.8550 0.6800 3.9750 2.1500 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0850 0.6800 5.2050 2.1200 ;
        RECT  4.9450 0.9400 5.2050 1.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.6650 -0.1800 4.7850 0.7300 ;
        RECT  3.4350 -0.1800 3.5550 0.7300 ;
        RECT  1.8600 -0.1800 1.9800 0.6400 ;
        RECT  0.5800 -0.1800 0.7000 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.6650 1.4700 4.7850 2.7900 ;
        RECT  3.4350 1.5000 3.5550 2.7900 ;
        RECT  2.0600 2.2300 2.1800 2.7900 ;
        RECT  0.6200 1.8800 0.7400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.9650 1.3300 4.3650 1.3300 4.3650 2.1200 4.2450 2.1200 4.2450 0.6800 4.3650 0.6800
                 4.3650 1.2100 4.9650 1.2100 ;
        POLYGON  3.7050 1.2400 3.5850 1.2400 3.5850 0.9700 3.1950 0.9700 3.1950 0.5600 2.5200 0.5600
                 2.5200 1.6300 2.6600 1.6300 2.6600 1.8700 2.5400 1.8700 2.5400 1.7500 2.4000 1.7500
                 2.4000 1.3500 2.0400 1.3500 2.0400 1.4700 1.9200 1.4700 1.9200 1.2300 2.4000 1.2300
                 2.4000 0.6400 2.2800 0.6400 2.2800 0.4000 2.4000 0.4000 2.4000 0.4400 3.3150 0.4400
                 3.3150 0.8500 3.7050 0.8500 ;
        POLYGON  3.0750 2.1100 1.7500 2.1100 1.7500 2.1500 1.1200 2.1500 1.1200 1.4300 1.3800 1.4300
                 1.3800 0.9000 0.3600 0.9000 0.3600 0.7800 1.5000 0.7800 1.5000 1.3100 1.5600 1.3100
                 1.5600 1.5500 1.2400 1.5500 1.2400 2.0300 1.6300 2.0300 1.6300 1.9900 2.9550 1.9900
                 2.9550 0.6800 3.0750 0.6800 ;
        POLYGON  2.2800 1.0600 1.8000 1.0600 1.8000 1.7900 1.4800 1.7900 1.4800 1.9100 1.3600 1.9100
                 1.3600 1.6700 1.6800 1.6700 1.6800 1.0600 1.6200 1.0600 1.6200 0.6400 1.2200 0.6400
                 1.2200 0.4000 1.3400 0.4000 1.3400 0.5200 1.7400 0.5200 1.7400 0.9400 2.1600 0.9400
                 2.1600 0.8200 2.2800 0.8200 ;
        POLYGON  1.2600 1.2200 1.0000 1.2200 1.0000 1.7600 0.2600 1.7600 0.2600 1.8800 0.1400 1.8800
                 0.1400 1.7600 0.1200 1.7600 0.1200 0.5200 0.1600 0.5200 0.1600 0.4000 0.2800 0.4000
                 0.2800 0.6400 0.2400 0.6400 0.2400 1.6400 0.8800 1.6400 0.8800 1.1000 1.2600 1.1000 ;
    END
END TLATNX1

MACRO TLATNTSCAX8
    CLASS CORE ;
    FOREIGN TLATNTSCAX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 0.8250 0.5650 1.0900 ;
        RECT  0.3250 0.7800 0.5650 1.0900 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9250 0.7600 1.0900 1.2300 ;
        RECT  0.9250 0.7600 1.0450 1.2600 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 0.8000 1.3850 1.2600 ;
        RECT  1.2300 0.7600 1.3800 1.1950 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3000 1.2250 9.4200 2.2050 ;
        RECT  9.2600 0.6450 9.3800 1.3450 ;
        RECT  6.7400 1.2250 9.4200 1.3450 ;
        RECT  7.6400 0.7650 9.3800 0.8850 ;
        RECT  8.3600 0.7150 8.6000 0.8850 ;
        RECT  8.4600 1.2250 8.5800 2.2050 ;
        RECT  7.5200 0.7150 7.7600 0.8350 ;
        RECT  7.6200 1.2250 7.7400 2.2100 ;
        RECT  6.7800 0.7750 6.9000 2.2100 ;
        RECT  6.7400 0.6550 6.8600 0.8950 ;
        RECT  6.7400 1.1750 6.9000 1.4350 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.8400 -0.1800 8.9600 0.6450 ;
        RECT  8.0000 -0.1800 8.1200 0.6450 ;
        RECT  7.1600 -0.1800 7.2800 0.6450 ;
        RECT  6.3200 -0.1800 6.4400 0.6400 ;
        RECT  5.0400 -0.1800 5.1600 0.7400 ;
        RECT  3.3500 0.4100 3.5900 0.5300 ;
        RECT  3.4700 -0.1800 3.5900 0.5300 ;
        RECT  1.0800 -0.1800 1.2000 0.6400 ;
        RECT  0.2400 -0.1800 0.3600 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.8800 1.4650 9.0000 2.7900 ;
        RECT  8.0400 1.4650 8.1600 2.7900 ;
        RECT  7.2000 1.4650 7.3200 2.7900 ;
        RECT  6.3600 1.7700 6.4800 2.7900 ;
        RECT  5.5200 1.7700 5.6400 2.7900 ;
        RECT  4.6600 1.6900 4.7800 2.7900 ;
        RECT  3.2500 2.0000 3.3700 2.7900 ;
        RECT  3.1300 2.0000 3.3700 2.1200 ;
        RECT  0.9600 1.6200 1.0800 2.7900 ;
        RECT  0.8400 1.6200 1.0800 1.7400 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.6200 1.2150 6.4000 1.2150 6.4000 1.6500 6.0600 1.6500 6.0600 2.2100 5.9400 2.2100
                 5.9400 1.6500 5.2200 1.6500 5.2200 2.2100 5.1000 2.2100 5.1000 1.5300 6.2800 1.5300
                 6.2800 1.0500 5.7600 1.0500 5.7600 0.8100 5.6800 0.8100 5.6800 0.5700 5.8000 0.5700
                 5.8000 0.6900 5.8800 0.6900 5.8800 0.9300 6.6200 0.9300 ;
        POLYGON  6.1600 1.4100 5.0400 1.4100 5.0400 1.2500 4.3000 1.2500 4.3000 2.0100 4.1800 2.0100
                 4.1800 1.4000 3.1300 1.4000 3.1300 1.2800 4.1800 1.2800 4.1800 1.1300 4.5600 1.1300
                 4.5600 0.6000 4.6800 0.6000 4.6800 1.1300 5.1600 1.1300 5.1600 1.2900 6.0400 1.2900
                 6.0400 1.1700 6.1600 1.1700 ;
        POLYGON  5.6400 1.1700 5.5200 1.1700 5.5200 1.0500 5.4400 1.0500 5.4400 0.9800 4.8000 0.9800
                 4.8000 0.4800 4.1900 0.4800 4.1900 0.7600 4.0700 0.7600 4.0700 1.0100 4.0600 1.0100
                 4.0600 1.1600 3.0100 1.1600 3.0100 1.5200 3.8500 1.5200 3.8500 1.8800 3.9700 1.8800
                 3.9700 2.0000 3.7300 2.0000 3.7300 1.6400 2.8900 1.6400 2.8900 1.3000 2.8500 1.3000
                 2.8500 1.0400 3.9400 1.0400 3.9400 0.8900 3.9500 0.8900 3.9500 0.6400 4.0700 0.6400
                 4.0700 0.3600 4.9200 0.3600 4.9200 0.8600 5.5600 0.8600 5.5600 0.9300 5.6400 0.9300 ;
        POLYGON  4.5400 2.2500 3.4900 2.2500 3.4900 1.8800 2.6700 1.8800 2.6700 2.0600 2.5500 2.0600
                 2.5500 1.9400 2.3700 1.9400 2.3700 0.8200 2.2500 0.8200 2.2500 0.7000 2.4900 0.7000
                 2.4900 1.7600 3.6100 1.7600 3.6100 2.1300 4.4200 2.1300 4.4200 1.3700 4.5400 1.3700 ;
        POLYGON  3.9500 0.4800 3.8300 0.4800 3.8300 0.7700 2.7300 0.7700 2.7300 1.6400 2.6100 1.6400
                 2.6100 0.5800 2.3450 0.5800 2.3450 0.5200 1.6250 0.5200 1.6250 1.5000 1.6800 1.5000
                 1.6800 1.6200 1.4400 1.6200 1.4400 1.5000 1.5050 1.5000 1.5050 0.6400 1.5000 0.6400
                 1.5000 0.4000 2.1100 0.4000 2.1100 0.3800 2.3500 0.3800 2.3500 0.4000 2.4650 0.4000
                 2.4650 0.4600 2.7300 0.4600 2.7300 0.6500 3.7100 0.6500 3.7100 0.3600 3.9500 0.3600 ;
        POLYGON  2.2500 2.0600 2.1300 2.0600 2.1300 1.9400 1.2000 1.9400 1.2000 1.5000 0.3800 1.5000
                 0.3800 1.6800 0.2600 1.6800 0.2600 1.3800 0.6850 1.3800 0.6850 0.6600 0.6600 0.6600
                 0.6600 0.4000 0.7800 0.4000 0.7800 0.5400 0.8050 0.5400 0.8050 1.3800 1.3200 1.3800
                 1.3200 1.8200 1.8900 1.8200 1.8900 0.6400 2.0100 0.6400 2.0100 1.8200 2.2500 1.8200 ;
    END
END TLATNTSCAX8

MACRO TLATNTSCAX6
    CLASS CORE ;
    FOREIGN TLATNTSCAX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 0.8200 0.5650 1.0900 ;
        RECT  0.3250 0.7600 0.5650 1.0900 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9250 0.7600 1.0900 1.2050 ;
        RECT  0.9250 0.7600 1.0450 1.2300 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 0.7600 1.3850 1.2500 ;
        RECT  1.2300 0.7600 1.3850 1.2200 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1924  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4450 1.1900 8.5650 2.2100 ;
        RECT  8.4450 0.4050 8.5650 1.0400 ;
        RECT  6.7400 1.1900 8.5650 1.3100 ;
        RECT  8.2650 0.9200 8.5650 1.0400 ;
        RECT  7.6050 1.0400 8.3850 1.3100 ;
        RECT  7.6050 0.4050 7.7250 2.2100 ;
        RECT  6.7400 1.1750 6.8900 1.4350 ;
        RECT  6.7650 0.4050 6.8850 2.2100 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  8.0250 -0.1800 8.1450 0.9200 ;
        RECT  7.1850 -0.1800 7.3050 0.9200 ;
        RECT  6.3450 -0.1800 6.4650 0.8300 ;
        RECT  4.9450 -0.1800 5.1850 0.3200 ;
        RECT  3.3550 -0.1800 3.5950 0.3400 ;
        RECT  1.0850 -0.1800 1.2050 0.6400 ;
        RECT  0.2450 -0.1800 0.3650 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  8.0250 1.4300 8.1450 2.7900 ;
        RECT  7.1850 1.4300 7.3050 2.7900 ;
        RECT  6.3450 1.7700 6.4650 2.7900 ;
        RECT  5.5050 1.7700 5.6250 2.7900 ;
        RECT  4.6650 1.5600 4.7850 2.7900 ;
        RECT  3.1950 2.1800 3.4350 2.3000 ;
        RECT  3.1950 2.1800 3.3150 2.7900 ;
        RECT  0.9650 1.6100 1.0850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.6050 1.2800 6.5050 1.2800 6.5050 1.6500 6.0450 1.6500 6.0450 2.2100 5.9250 2.2100
                 5.9250 1.6500 5.2050 1.6500 5.2050 2.2100 5.0850 2.2100 5.0850 1.5300 6.3850 1.5300
                 6.3850 1.1600 5.7850 1.1600 5.7850 0.8100 5.7050 0.8100 5.7050 0.5700 5.8250 0.5700
                 5.8250 0.6900 5.9050 0.6900 5.9050 1.0400 6.6050 1.0400 ;
        POLYGON  6.2650 1.4000 6.1450 1.4000 6.1450 1.4100 5.0250 1.4100 5.0250 1.1800 4.3050 1.1800
                 4.3050 1.5000 4.1850 1.5000 4.1850 1.6200 4.3050 1.6200 4.3050 2.0100 4.0650 2.0100
                 4.0650 1.5000 3.1750 1.5000 3.1750 1.3800 4.1850 1.3800 4.1850 1.0600 4.4650 1.0600
                 4.4650 0.6800 4.7050 0.6800 4.7050 0.8000 4.5850 0.8000 4.5850 1.0600 5.0250 1.0600
                 5.0250 1.0500 5.1450 1.0500 5.1450 1.2900 6.0250 1.2900 6.0250 1.2800 6.2650 1.2800 ;
        POLYGON  5.6650 1.1700 5.5450 1.1700 5.5450 1.0500 5.4650 1.0500 5.4650 0.9300 4.9350 0.9300
                 4.9350 0.5600 4.2150 0.5600 4.2150 0.8000 4.0750 0.8000 4.0750 0.9200 4.0650 0.9200
                 4.0650 1.1800 3.0550 1.1800 3.0550 1.6200 3.7950 1.6200 3.7950 1.7000 3.9150 1.7000
                 3.9150 1.8200 3.6750 1.8200 3.6750 1.7400 2.9350 1.7400 2.9350 1.1800 2.8550 1.1800
                 2.8550 1.0600 3.9450 1.0600 3.9450 0.8000 3.9550 0.8000 3.9550 0.6800 4.0950 0.6800
                 4.0950 0.4400 5.0550 0.4400 5.0550 0.8100 5.5850 0.8100 5.5850 0.9300 5.6650 0.9300 ;
        POLYGON  4.6650 1.4200 4.5450 1.4200 4.5450 2.2500 3.6150 2.2500 3.6150 2.0600 2.5550 2.0600
                 2.5550 1.8200 2.3750 1.8200 2.3750 0.8600 2.2550 0.8600 2.2550 0.7400 2.4950 0.7400
                 2.4950 1.7000 2.6750 1.7000 2.6750 1.9400 3.7350 1.9400 3.7350 2.1300 4.4250 2.1300
                 4.4250 1.3000 4.6650 1.3000 ;
        POLYGON  3.9750 0.5200 3.8350 0.5200 3.8350 0.5800 2.7350 0.5800 2.7350 1.3000 2.8150 1.3000
                 2.8150 1.5600 2.6950 1.5600 2.6950 1.4200 2.6150 1.4200 2.6150 0.5800 2.5000 0.5800
                 2.5000 0.5400 1.6250 0.5400 1.6250 1.5500 1.6850 1.5500 1.6850 1.6700 1.4450 1.6700
                 1.4450 1.5500 1.5050 1.5500 1.5050 0.4000 1.6250 0.4000 1.6250 0.4200 2.6200 0.4200
                 2.6200 0.4600 3.7150 0.4600 3.7150 0.4000 3.9750 0.4000 ;
        POLYGON  2.2550 1.9100 1.2050 1.9100 1.2050 1.4900 0.5050 1.4900 0.5050 1.6700 0.2650 1.6700
                 0.2650 1.5500 0.3850 1.5500 0.3850 1.3700 0.6850 1.3700 0.6850 0.6400 0.6650 0.6400
                 0.6650 0.4000 0.7850 0.4000 0.7850 0.5200 0.8050 0.5200 0.8050 1.3700 1.3250 1.3700
                 1.3250 1.7900 2.0150 1.7900 2.0150 0.9200 1.8950 0.9200 1.8950 0.6800 2.0150 0.6800
                 2.0150 0.8000 2.1350 0.8000 2.1350 1.6400 2.2550 1.6400 ;
    END
END TLATNTSCAX6

MACRO TLATNTSCAX4
    CLASS CORE ;
    FOREIGN TLATNTSCAX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7050 0.5900 6.8250 2.2100 ;
        RECT  5.8700 1.0250 6.8250 1.1450 ;
        RECT  5.8650 0.8850 6.0200 1.0250 ;
        RECT  5.8850 0.8850 6.0050 1.6800 ;
        RECT  5.8650 1.5600 5.9850 2.2100 ;
        RECT  5.8650 0.5900 5.9850 1.0250 ;
        END
    END ECK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.4350 1.2950 ;
        RECT  0.3150 1.0550 0.4350 1.2950 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1650 1.1450 1.4000 ;
        RECT  0.7950 1.1650 1.1450 1.3750 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1350 1.5200 1.4350 1.7550 ;
        END
    END CK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  7.1250 -0.1800 7.2450 0.6400 ;
        RECT  6.2850 -0.1800 6.4050 0.6400 ;
        RECT  5.4450 -0.1800 5.5650 0.6400 ;
        RECT  4.4150 -0.1800 4.5350 0.9000 ;
        RECT  3.0650 0.6800 3.3050 0.8000 ;
        RECT  3.1850 -0.1800 3.3050 0.8000 ;
        RECT  0.9550 0.6850 1.1950 0.8050 ;
        RECT  0.9550 -0.1800 1.0750 0.8050 ;
        RECT  0.1750 -0.1800 0.2950 0.8650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  7.1250 1.5600 7.2450 2.7900 ;
        RECT  6.2850 1.5600 6.4050 2.7900 ;
        RECT  5.4450 1.6000 5.5650 2.7900 ;
        RECT  4.6250 1.8000 4.7450 2.7900 ;
        RECT  4.6050 1.5600 4.7250 1.9200 ;
        RECT  3.2550 2.2900 3.4950 2.7900 ;
        RECT  1.0150 1.9000 1.1350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7650 1.3850 5.4450 1.3850 5.4450 1.4800 5.1450 1.4800 5.1450 2.2100 5.0250 2.2100
                 5.0250 1.3600 5.3250 1.3600 5.3250 0.8800 5.0550 0.8800 5.0550 0.6400 5.1750 0.6400
                 5.1750 0.7600 5.4450 0.7600 5.4450 1.2650 5.7650 1.2650 ;
        POLYGON  5.2050 1.2400 5.0850 1.2400 5.0850 1.1400 4.1750 1.1400 4.1750 0.5400 3.7650 0.5400
                 3.7650 0.7400 3.8150 0.7400 3.8150 1.5700 3.9750 1.5700 3.9750 1.6900 3.6950 1.6900
                 3.6950 1.0400 2.8250 1.0400 2.8250 0.5600 2.3050 0.5600 2.3050 1.6400 2.1850 1.6400
                 2.1850 0.4400 2.5650 0.4400 2.5650 0.3600 2.8050 0.3600 2.8050 0.4400 2.9450 0.4400
                 2.9450 0.9200 3.5450 0.9200 3.5450 0.6200 3.6450 0.6200 3.6450 0.4200 4.2950 0.4200
                 4.2950 1.0200 5.0850 1.0200 5.0850 1.0000 5.2050 1.0000 ;
        POLYGON  4.8650 1.4200 4.3050 1.4200 4.3050 1.9300 3.1450 1.9300 3.1450 1.6000 3.0250 1.6000
                 3.0250 1.4800 3.2650 1.4800 3.2650 1.8100 4.1850 1.8100 4.1850 1.3800 3.9350 1.3800
                 3.9350 0.6600 4.0550 0.6600 4.0550 1.2600 4.3050 1.2600 4.3050 1.3000 4.8650 1.3000 ;
        POLYGON  4.5050 2.1800 4.0000 2.1800 4.0000 2.1700 2.4250 2.1700 2.4250 0.6800 2.6650 0.6800
                 2.6650 0.8000 2.5450 0.8000 2.5450 1.8600 2.7050 1.8600 2.7050 2.0500 4.1200 2.0500
                 4.1200 2.0600 4.5050 2.0600 ;
        POLYGON  3.4850 1.2800 3.3650 1.2800 3.3650 1.3400 2.6650 1.3400 2.6650 1.2200 3.2450 1.2200
                 3.2450 1.1600 3.4850 1.1600 ;
        POLYGON  2.2850 2.0000 2.1650 2.0000 2.1650 1.8800 1.9450 1.8800 1.9450 0.5050 1.4350 0.5050
                 1.4350 1.0450 0.6750 1.0450 0.6750 1.9600 0.3150 1.9600 0.3150 1.8400 0.5550 1.8400
                 0.5550 0.8050 0.5950 0.8050 0.5950 0.6250 0.7150 0.6250 0.7150 0.9250 1.3150 0.9250
                 1.3150 0.3850 2.0650 0.3850 2.0650 1.7600 2.2850 1.7600 ;
        POLYGON  1.8250 1.4000 1.6750 1.4000 1.6750 1.9950 1.5550 1.9950 1.5550 2.1150 1.4350 2.1150
                 1.4350 1.8750 1.5550 1.8750 1.5550 0.6250 1.6750 0.6250 1.6750 1.1600 1.8250 1.1600 ;
    END
END TLATNTSCAX4

MACRO TLATNTSCAX3
    CLASS CORE ;
    FOREIGN TLATNTSCAX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.2500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 0.8200 0.5650 1.0900 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 0.7600 1.0900 1.1800 ;
        RECT  0.9250 0.8000 1.0450 1.2400 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 0.7600 1.3850 1.2400 ;
        RECT  1.2300 0.7600 1.3850 1.2150 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9950 0.5900 7.1150 0.8300 ;
        RECT  6.8150 0.7100 7.1150 0.8300 ;
        RECT  6.8250 1.3100 6.9450 2.2000 ;
        RECT  6.1600 0.8300 6.9350 0.9500 ;
        RECT  6.1600 1.3100 6.9450 1.4300 ;
        RECT  6.1600 0.8300 6.3100 1.1450 ;
        RECT  5.9850 1.4300 6.2800 1.5500 ;
        RECT  6.1600 0.7100 6.2800 1.5500 ;
        RECT  6.1550 0.5900 6.2750 0.8300 ;
        RECT  5.9850 1.4300 6.1050 2.2000 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.2500 0.1800 ;
        RECT  6.5750 -0.1800 6.6950 0.6400 ;
        RECT  5.6750 -0.1800 5.7950 0.5300 ;
        RECT  4.6050 -0.1800 4.8450 0.3800 ;
        RECT  3.1950 0.7000 3.4350 0.8200 ;
        RECT  3.2350 -0.1800 3.3550 0.8200 ;
        RECT  0.9850 -0.1800 1.1050 0.6400 ;
        RECT  0.1450 -0.1800 0.2650 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.2500 2.7900 ;
        RECT  6.4050 1.5500 6.5250 2.7900 ;
        RECT  5.5650 1.6400 5.6850 2.7900 ;
        RECT  4.7250 1.5500 4.8450 2.7900 ;
        RECT  3.0350 2.1400 3.2750 2.2600 ;
        RECT  3.0350 2.1400 3.1550 2.7900 ;
        RECT  0.9450 1.6000 1.0650 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.0400 1.1900 5.5650 1.1900 5.5650 1.5200 5.2650 1.5200 5.2650 2.2000 5.1450 2.2000
                 5.1450 1.4000 5.4450 1.4000 5.4450 0.9200 5.3650 0.9200 5.3650 0.6800 5.4850 0.6800
                 5.4850 0.8000 5.5650 0.8000 5.5650 1.0700 6.0400 1.0700 ;
        POLYGON  5.3250 1.2800 5.1250 1.2800 5.1250 0.6200 3.9550 0.6200 3.9550 0.7600 3.9150 0.7600
                 3.9150 1.3000 2.9550 1.3000 2.9550 1.6600 3.7550 1.6600 3.7550 1.8900 3.8750 1.8900
                 3.8750 2.0100 3.6350 2.0100 3.6350 1.7800 2.8350 1.7800 2.8350 1.3000 2.6950 1.3000
                 2.6950 1.1800 3.7950 1.1800 3.7950 0.6400 3.8350 0.6400 3.8350 0.5000 5.2450 0.5000
                 5.2450 1.0400 5.3250 1.0400 ;
        POLYGON  5.0050 1.2600 4.3650 1.2600 4.3650 1.6100 4.4850 1.6100 4.4850 1.7300 4.2450 1.7300
                 4.2450 1.5400 3.0750 1.5400 3.0750 1.4200 4.2450 1.4200 4.2450 0.8600 4.1250 0.8600
                 4.1250 0.7400 4.3650 0.7400 4.3650 1.1400 5.0050 1.1400 ;
        POLYGON  4.5850 2.2500 3.3950 2.2500 3.3950 2.0200 2.5150 2.0200 2.5150 2.0700 2.3950 2.0700
                 2.3950 1.9500 2.2150 1.9500 2.2150 0.6400 2.3350 0.6400 2.3350 1.8300 2.5150 1.8300
                 2.5150 1.9000 3.5150 1.9000 3.5150 2.1300 4.4650 2.1300 4.4650 2.0100 4.5850 2.0100 ;
        POLYGON  3.7150 0.4800 3.6750 0.4800 3.6750 1.0600 2.9550 1.0600 2.9550 0.5200 2.5750 0.5200
                 2.5750 1.5700 2.7150 1.5700 2.7150 1.6900 2.4550 1.6900 2.4550 0.5200 1.6250 0.5200
                 1.6250 1.4800 1.5450 1.4800 1.5450 1.7200 1.4250 1.7200 1.4250 1.3600 1.5050 1.3600
                 1.5050 0.6400 1.4050 0.6400 1.4050 0.4000 1.9950 0.4000 1.9950 0.3600 2.2350 0.3600
                 2.2350 0.4000 3.0750 0.4000 3.0750 0.9400 3.5550 0.9400 3.5550 0.4800 3.4750 0.4800
                 3.4750 0.3600 3.7150 0.3600 ;
        POLYGON  2.0950 2.0700 1.9750 2.0700 1.9750 1.9600 1.1850 1.9600 1.1850 1.4800 0.4250 1.4800
                 0.4250 1.7200 0.3050 1.7200 0.3050 1.3600 0.6850 1.3600 0.6850 0.7000 0.5650 0.7000
                 0.5650 0.4000 0.6850 0.4000 0.6850 0.5800 0.8050 0.5800 0.8050 1.3600 1.3050 1.3600
                 1.3050 1.8400 1.9750 1.8400 1.9750 0.8800 1.7950 0.8800 1.7950 0.6400 1.9150 0.6400
                 1.9150 0.7600 2.0950 0.7600 ;
    END
END TLATNTSCAX3

MACRO TLATNTSCAX20
    CLASS CORE ;
    FOREIGN TLATNTSCAX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 16.5300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 1.0400 0.2900 1.3350 ;
        RECT  0.0700 1.1300 0.2200 1.4350 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8200 1.0400 0.9400 1.2800 ;
        RECT  0.6800 1.1600 0.9400 1.2800 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2300 1.4350 1.3800 ;
        RECT  1.1800 1.1000 1.4200 1.3800 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.6080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  16.1000 1.2050 16.2200 2.2050 ;
        RECT  16.1000 0.4050 16.2200 1.0300 ;
        RECT  9.3500 1.2050 16.2200 1.3250 ;
        RECT  15.9200 0.9100 16.2200 1.0300 ;
        RECT  15.2600 1.0300 16.0400 1.3250 ;
        RECT  15.2600 0.4050 15.3800 2.2100 ;
        RECT  14.4200 0.4050 14.5400 2.2100 ;
        RECT  13.5800 1.0300 14.5400 1.3250 ;
        RECT  13.5800 0.4050 13.7000 2.2100 ;
        RECT  12.7400 0.4050 12.8600 2.2100 ;
        RECT  11.9000 1.0300 12.8600 1.3250 ;
        RECT  11.9000 0.4050 12.0200 2.2100 ;
        RECT  11.0600 1.2050 11.1800 2.2100 ;
        RECT  10.8800 0.7900 11.1800 0.9100 ;
        RECT  11.0600 0.4050 11.1800 0.9100 ;
        RECT  10.2200 1.0300 11.0000 1.3250 ;
        RECT  10.8800 0.7900 11.0000 1.3250 ;
        RECT  10.2200 0.4050 10.3400 2.2100 ;
        RECT  9.3800 0.4000 9.5000 2.2100 ;
        RECT  9.3500 1.1750 9.5000 1.4350 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 16.5300 0.1800 ;
        RECT  15.6800 -0.1800 15.8000 0.9100 ;
        RECT  14.8400 -0.1800 14.9600 0.9100 ;
        RECT  14.0000 -0.1800 14.1200 0.9100 ;
        RECT  13.1600 -0.1800 13.2800 0.9100 ;
        RECT  12.3200 -0.1800 12.4400 0.9100 ;
        RECT  11.4800 -0.1800 11.6000 0.9100 ;
        RECT  10.6400 -0.1800 10.7600 0.9100 ;
        RECT  9.8000 -0.1800 9.9200 0.9100 ;
        RECT  8.9600 -0.1800 9.0800 0.8700 ;
        RECT  7.6400 0.4600 7.8800 0.5800 ;
        RECT  7.6400 -0.1800 7.7600 0.5800 ;
        RECT  6.3600 0.4600 6.6000 0.5800 ;
        RECT  6.3600 -0.1800 6.4800 0.5800 ;
        RECT  5.1400 -0.1800 5.2600 0.6400 ;
        RECT  4.3000 -0.1800 4.4200 0.6400 ;
        RECT  2.9700 0.4700 3.2100 0.5900 ;
        RECT  2.9700 -0.1800 3.0900 0.5900 ;
        RECT  0.9800 -0.1800 1.2200 0.3400 ;
        RECT  0.1400 -0.1800 0.2600 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 16.5300 2.7900 ;
        RECT  15.6800 1.4450 15.8000 2.7900 ;
        RECT  14.8400 1.4450 14.9600 2.7900 ;
        RECT  14.0000 1.4450 14.1200 2.7900 ;
        RECT  13.1600 1.4450 13.2800 2.7900 ;
        RECT  12.3200 1.4450 12.4400 2.7900 ;
        RECT  11.4800 1.4450 11.6000 2.7900 ;
        RECT  10.6400 1.4450 10.7600 2.7900 ;
        RECT  9.8000 1.4450 9.9200 2.7900 ;
        RECT  8.9600 1.7100 9.0800 2.7900 ;
        RECT  8.1200 1.7100 8.2400 2.7900 ;
        RECT  7.2800 1.7100 7.4000 2.7900 ;
        RECT  6.4400 1.7100 6.5600 2.7900 ;
        RECT  5.6000 1.7100 5.7200 2.7900 ;
        RECT  4.7000 2.0300 4.9400 2.1500 ;
        RECT  4.7000 2.0300 4.8200 2.7900 ;
        RECT  3.7400 2.0600 3.9800 2.1800 ;
        RECT  3.7400 2.0600 3.8600 2.7900 ;
        RECT  3.0700 2.0300 3.1900 2.7900 ;
        RECT  0.9800 1.5000 1.1000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.2300 1.2300 9.0200 1.2300 9.0200 1.5900 8.6600 1.5900 8.6600 2.2100 8.5400 2.2100
                 8.5400 1.5900 7.8200 1.5900 7.8200 2.2100 7.7000 2.2100 7.7000 1.5900 6.9800 1.5900
                 6.9800 2.2100 6.8600 2.2100 6.8600 1.5900 6.1400 1.5900 6.1400 2.2100 6.0200 2.2100
                 6.0200 1.5900 5.3000 1.5900 5.3000 2.2100 5.1800 2.2100 5.1800 1.4700 8.9000 1.4700
                 8.9000 1.1100 8.3400 1.1100 8.3400 0.8200 5.8400 0.8200 5.8400 0.7700 5.7200 0.7700
                 5.7200 0.6500 5.9600 0.6500 5.9600 0.7000 7.0000 0.7000 7.0000 0.6500 7.2400 0.6500
                 7.2400 0.7000 8.3400 0.7000 8.3400 0.5900 8.4600 0.5900 8.4600 0.9900 9.0200 0.9900
                 9.0200 1.1100 9.2300 1.1100 ;
        POLYGON  8.7800 1.3500 5.0600 1.3500 5.0600 1.9100 3.7100 1.9100 3.7100 1.6700 2.6300 1.6700
                 2.6300 1.2900 2.5500 1.2900 2.5500 1.0500 2.6300 1.0500 2.6300 0.9500 3.5700 0.9500
                 3.5700 0.6000 3.8100 0.6000 3.8100 0.7200 3.6900 0.7200 3.6900 1.0700 2.7500 1.0700
                 2.7500 1.5500 3.8300 1.5500 3.8300 1.7900 4.9400 1.7900 4.9400 1.2300 8.7800 1.2300 ;
        POLYGON  8.0200 1.1100 4.8200 1.1100 4.8200 1.4300 4.3400 1.4300 4.3400 1.5500 4.4600 1.5500
                 4.4600 1.6700 4.2200 1.6700 4.2200 1.4300 2.8700 1.4300 2.8700 1.1900 2.9900 1.1900
                 2.9900 1.3100 4.7000 1.3100 4.7000 0.7100 4.7200 0.7100 4.7200 0.5900 4.8400 0.5900
                 4.8400 0.8300 4.8200 0.8300 4.8200 0.9900 8.0200 0.9900 ;
        POLYGON  4.5600 1.1900 4.0200 1.1900 4.0200 1.0700 4.4400 1.0700 4.4400 0.9500 4.0600 0.9500
                 4.0600 0.4800 3.4500 0.4800 3.4500 0.8300 2.4300 0.8300 2.4300 1.7900 2.5500 1.7900
                 2.5500 1.9100 2.3100 1.9100 2.3100 0.6100 2.3300 0.6100 2.3300 0.4900 2.4500 0.4900
                 2.4500 0.7100 3.3300 0.7100 3.3300 0.3600 4.1800 0.3600 4.1800 0.8300 4.5600 0.8300 ;
        POLYGON  3.5900 2.1100 3.3500 2.1100 3.3500 1.9100 2.9500 1.9100 2.9500 2.1500 2.7100 2.1500
                 2.7100 2.2500 2.4700 2.2500 2.4700 2.1500 2.0700 2.1500 2.0700 2.0900 1.5400 2.0900
                 1.5400 1.8600 1.4000 1.8600 1.4000 1.5000 1.5550 1.5000 1.5550 0.8600 1.4600 0.8600
                 1.4600 0.7400 1.7000 0.7400 1.7000 0.8600 1.6750 0.8600 1.6750 1.6200 1.5200 1.6200
                 1.5200 1.7400 1.6600 1.7400 1.6600 1.9700 2.0700 1.9700 2.0700 0.8500 2.1900 0.8500
                 2.1900 2.0300 2.8300 2.0300 2.8300 1.7900 3.4700 1.7900 3.4700 1.9900 3.5900 1.9900 ;
        POLYGON  2.0300 0.7300 1.9500 0.7300 1.9500 1.8500 1.8300 1.8500 1.8300 0.6200 1.2100 0.6200
                 1.2100 0.6800 0.6800 0.6800 0.6800 0.9200 0.5300 0.9200 0.5300 1.5750 0.4600 1.5750
                 0.4600 1.6950 0.3400 1.6950 0.3400 1.4550 0.4100 1.4550 0.4100 0.8000 0.5600 0.8000
                 0.5600 0.5600 1.0900 0.5600 1.0900 0.5000 1.9100 0.5000 1.9100 0.4900 2.0300 0.4900 ;
    END
END TLATNTSCAX20

MACRO TLATNTSCAX2
    CLASS CORE ;
    FOREIGN TLATNTSCAX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3250 0.8200 0.5650 1.2200 ;
        RECT  0.3050 0.8200 0.5650 1.0900 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 0.7600 1.0900 1.1750 ;
        RECT  0.9250 0.8100 1.0450 1.2450 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.7600 1.3800 1.2200 ;
        RECT  1.2450 0.7600 1.3650 1.2450 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9950 0.5900 6.1150 0.8300 ;
        RECT  5.8700 0.7100 6.0200 1.1450 ;
        RECT  5.8650 1.1450 5.9900 1.2650 ;
        RECT  5.8650 1.1450 5.9850 1.9900 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  6.4150 -0.1800 6.5350 0.6400 ;
        RECT  5.5150 -0.1800 5.6350 0.5300 ;
        RECT  4.6550 -0.1800 4.7750 0.4000 ;
        RECT  3.1850 0.7000 3.4250 0.8200 ;
        RECT  3.2250 -0.1800 3.3450 0.8200 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  6.2850 1.3400 6.4050 2.7900 ;
        RECT  5.4450 1.3600 5.5650 2.7900 ;
        RECT  4.6050 1.4800 4.7250 2.7900 ;
        RECT  3.0250 2.1400 3.2650 2.2600 ;
        RECT  3.0250 2.1400 3.1450 2.7900 ;
        RECT  0.9250 1.6050 1.0450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7450 1.1800 5.1850 1.1800 5.1850 1.4400 5.1450 1.4400 5.1450 1.6000 5.0250 1.6000
                 5.0250 1.3200 5.0650 1.3200 5.0650 1.0600 5.3050 1.0600 5.3050 0.8600 5.1850 0.8600
                 5.1850 0.7400 5.4250 0.7400 5.4250 1.0600 5.7450 1.0600 ;
        POLYGON  5.2650 0.5200 5.0650 0.5200 5.0650 0.6400 4.4150 0.6400 4.4150 0.5600 3.9450 0.5600
                 3.9450 0.7600 3.9050 0.7600 3.9050 1.3000 2.9450 1.3000 2.9450 1.6600 3.7450 1.6600
                 3.7450 1.8900 3.8650 1.8900 3.8650 2.0100 3.6250 2.0100 3.6250 1.7800 2.8250 1.7800
                 2.8250 1.3000 2.6850 1.3000 2.6850 1.1800 3.7850 1.1800 3.7850 0.6400 3.8250 0.6400
                 3.8250 0.4400 4.5350 0.4400 4.5350 0.5200 4.9450 0.5200 4.9450 0.4000 5.2650 0.4000 ;
        POLYGON  4.9450 1.2000 4.2950 1.2000 4.2950 1.4200 4.3050 1.4200 4.3050 1.6600 4.1850 1.6600
                 4.1850 1.5400 3.0650 1.5400 3.0650 1.4200 4.1750 1.4200 4.1750 0.6800 4.2950 0.6800
                 4.2950 1.0800 4.9450 1.0800 ;
        POLYGON  4.4650 2.2500 3.3850 2.2500 3.3850 2.0200 2.5050 2.0200 2.5050 2.0700 2.3850 2.0700
                 2.3850 1.9500 2.2050 1.9500 2.2050 0.6400 2.3250 0.6400 2.3250 1.8300 2.5050 1.8300
                 2.5050 1.9000 3.5050 1.9000 3.5050 2.1300 4.3450 2.1300 4.3450 1.8200 4.4650 1.8200 ;
        POLYGON  3.7050 0.4800 3.6650 0.4800 3.6650 1.0600 2.9450 1.0600 2.9450 0.5200 2.5650 0.5200
                 2.5650 1.5700 2.7050 1.5700 2.7050 1.6900 2.4450 1.6900 2.4450 0.5200 1.6200 0.5200
                 1.6200 1.6050 1.5250 1.6050 1.5250 1.7250 1.4050 1.7250 1.4050 1.4850 1.5000 1.4850
                 1.5000 0.6400 1.3950 0.6400 1.3950 0.4000 1.9850 0.4000 1.9850 0.3600 2.2250 0.3600
                 2.2250 0.4000 3.0650 0.4000 3.0650 0.9400 3.5450 0.9400 3.5450 0.4800 3.4650 0.4800
                 3.4650 0.3600 3.7050 0.3600 ;
        POLYGON  2.0850 2.0700 1.9650 2.0700 1.9650 1.9650 1.1650 1.9650 1.1650 1.4850 0.4050 1.4850
                 0.4050 1.7250 0.2850 1.7250 0.2850 1.3650 0.6850 1.3650 0.6850 0.7000 0.5550 0.7000
                 0.5550 0.4000 0.6750 0.4000 0.6750 0.5800 0.8050 0.5800 0.8050 1.3650 1.2850 1.3650
                 1.2850 1.8450 1.9650 1.8450 1.9650 0.8800 1.7850 0.8800 1.7850 0.6400 1.9050 0.6400
                 1.9050 0.7600 2.0850 0.7600 ;
    END
END TLATNTSCAX2

MACRO TLATNTSCAX16
    CLASS CORE ;
    FOREIGN TLATNTSCAX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.2100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 0.8450 0.5650 1.1000 ;
        RECT  0.2650 0.9800 0.5050 1.2100 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9250 0.7600 1.0900 1.2050 ;
        RECT  0.9250 0.7600 1.0450 1.2300 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 0.7600 1.3850 1.2500 ;
        RECT  1.2300 0.7600 1.3850 1.2200 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.5350 1.3450 13.6550 2.2050 ;
        RECT  8.4800 1.2250 13.5550 1.3450 ;
        RECT  13.4350 0.6550 13.5550 1.4650 ;
        RECT  12.6550 0.7750 13.5550 0.8950 ;
        RECT  12.6950 1.2250 12.8150 2.2050 ;
        RECT  12.5350 0.7250 12.7750 0.8450 ;
        RECT  11.8550 1.2250 11.9750 2.2050 ;
        RECT  11.7550 0.6550 11.8750 1.3450 ;
        RECT  10.9750 0.7750 11.8750 0.8950 ;
        RECT  11.0150 1.2250 11.1350 2.2100 ;
        RECT  10.8550 0.7250 11.0950 0.8450 ;
        RECT  10.1750 1.2250 10.2950 2.2100 ;
        RECT  10.0750 0.6550 10.1950 1.3450 ;
        RECT  9.2950 0.7750 10.1950 0.8950 ;
        RECT  9.3350 1.2250 9.4550 2.2100 ;
        RECT  9.1750 0.7250 9.4150 0.8450 ;
        RECT  8.4800 1.1750 8.6300 1.4350 ;
        RECT  8.4950 0.7850 8.6150 2.2100 ;
        RECT  8.3950 0.6650 8.5150 0.9050 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.2100 0.1800 ;
        RECT  13.8550 -0.1800 13.9750 0.6550 ;
        RECT  13.0150 -0.1800 13.1350 0.6550 ;
        RECT  12.1750 -0.1800 12.2950 0.6550 ;
        RECT  11.3350 -0.1800 11.4550 0.6550 ;
        RECT  10.4950 -0.1800 10.6150 0.6550 ;
        RECT  9.6550 -0.1800 9.7750 0.6550 ;
        RECT  8.8150 -0.1800 8.9350 0.6500 ;
        RECT  7.9750 -0.1800 8.0950 0.6500 ;
        RECT  6.4550 0.4700 6.6950 0.5900 ;
        RECT  6.4550 -0.1800 6.5750 0.5900 ;
        RECT  5.2350 -0.1800 5.3550 0.7600 ;
        RECT  4.1550 -0.1800 4.3950 0.3200 ;
        RECT  3.1950 0.4100 3.4350 0.5300 ;
        RECT  3.3150 -0.1800 3.4350 0.5300 ;
        RECT  1.0050 -0.1800 1.1250 0.6400 ;
        RECT  0.1650 -0.1800 0.2850 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.2100 2.7900 ;
        RECT  13.9550 1.4650 14.0750 2.7900 ;
        RECT  13.1150 1.4650 13.2350 2.7900 ;
        RECT  12.2750 1.4650 12.3950 2.7900 ;
        RECT  11.4350 1.4650 11.5550 2.7900 ;
        RECT  10.5950 1.4650 10.7150 2.7900 ;
        RECT  9.7550 1.4650 9.8750 2.7900 ;
        RECT  8.9150 1.4650 9.0350 2.7900 ;
        RECT  8.0750 1.7200 8.1950 2.7900 ;
        RECT  7.2350 1.7200 7.3550 2.7900 ;
        RECT  6.3950 1.7200 6.5150 2.7900 ;
        RECT  5.5550 1.7200 5.6750 2.7900 ;
        RECT  4.7150 1.6900 4.8350 2.7900 ;
        RECT  3.8150 2.2300 3.9350 2.7900 ;
        RECT  2.7650 1.9800 3.0050 2.1000 ;
        RECT  2.7650 1.9800 2.8850 2.7900 ;
        RECT  0.8850 1.6100 1.0050 2.7900 ;
        RECT  0.7650 1.6100 1.0050 1.7300 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2750 1.2400 8.1350 1.2400 8.1350 1.6000 7.7750 1.6000 7.7750 2.2100 7.6550 2.2100
                 7.6550 1.6000 6.9350 1.6000 6.9350 2.2100 6.8150 2.2100 6.8150 1.6000 6.0950 1.6000
                 6.0950 2.2100 5.9750 2.2100 5.9750 1.6000 5.2550 1.6000 5.2550 2.2100 5.1350 2.2100
                 5.1350 1.4800 8.0150 1.4800 8.0150 1.1200 7.3750 1.1200 7.3750 0.8400 7.2350 0.8400
                 7.2350 0.8300 5.9350 0.8300 5.9350 0.7800 5.8150 0.7800 5.8150 0.6600 6.0550 0.6600
                 6.0550 0.7100 7.2350 0.7100 7.2350 0.6000 7.3550 0.6000 7.3550 0.7200 7.4950 0.7200
                 7.4950 1.0000 8.2750 1.0000 ;
        POLYGON  7.8950 1.3600 4.5950 1.3600 4.5950 1.8100 4.4150 1.8100 4.4150 2.2100 4.2950 2.2100
                 4.2950 1.6900 4.4750 1.6900 4.4750 1.3100 3.1550 1.3100 3.1550 1.3700 3.0350 1.3700
                 3.0350 1.1300 3.1550 1.1300 3.1550 1.1900 4.6350 1.1900 4.6350 0.6800 4.8750 0.6800
                 4.8750 0.8000 4.7550 0.8000 4.7550 1.2400 7.8950 1.2400 ;
        POLYGON  7.2550 1.1200 5.5750 1.1200 5.5750 1.0000 4.9950 1.0000 4.9950 0.5600 4.5150 0.5600
                 4.5150 0.6400 4.0350 0.6400 4.0350 0.7600 3.9150 0.7600 3.9150 1.0100 2.9150 1.0100
                 2.9150 1.4900 3.4850 1.4900 3.4850 1.7500 3.6050 1.7500 3.6050 1.8700 3.3650 1.8700
                 3.3650 1.6100 2.7950 1.6100 2.7950 1.2600 2.7150 1.2600 2.7150 0.8900 3.7950 0.8900
                 3.7950 0.6400 3.9150 0.6400 3.9150 0.5200 4.3950 0.5200 4.3950 0.4400 5.1150 0.4400
                 5.1150 0.8800 5.6950 0.8800 5.6950 1.0000 7.2550 1.0000 ;
        POLYGON  4.3550 1.5500 4.1750 1.5500 4.1750 2.1100 3.1250 2.1100 3.1250 1.8600 2.6450 1.8600
                 2.6450 1.9200 2.3050 1.9200 2.3050 2.0400 2.1850 2.0400 2.1850 1.9200 2.1050 1.9200
                 2.1050 0.7400 2.2350 0.7400 2.2350 0.6200 2.3550 0.6200 2.3550 0.8600 2.2250 0.8600
                 2.2250 1.8000 2.5250 1.8000 2.5250 1.7400 3.2450 1.7400 3.2450 1.9900 4.0550 1.9900
                 4.0550 1.4300 4.3550 1.4300 ;
        POLYGON  3.7950 0.4800 3.6750 0.4800 3.6750 0.7700 2.9550 0.7700 2.9550 0.5000 2.5950 0.5000
                 2.5950 1.1000 2.4650 1.1000 2.4650 1.6200 2.3450 1.6200 2.3450 0.9800 2.4750 0.9800
                 2.4750 0.5000 1.6250 0.5000 1.6250 1.6100 1.3650 1.6100 1.3650 1.4900 1.5050 1.4900
                 1.5050 0.6400 1.4250 0.6400 1.4250 0.3800 2.0350 0.3800 2.0350 0.3600 2.2750 0.3600
                 2.2750 0.3800 3.0750 0.3800 3.0750 0.6500 3.5550 0.6500 3.5550 0.3600 3.7950 0.3600 ;
        POLYGON  1.9350 1.9400 1.8850 1.9400 1.8850 2.0600 1.7650 2.0600 1.7650 1.9400 1.1250 1.9400
                 1.1250 1.4900 0.3050 1.4900 0.3050 1.6700 0.1850 1.6700 0.1850 1.3700 0.6850 1.3700
                 0.6850 0.7250 0.5850 0.7250 0.5850 0.4000 0.7050 0.4000 0.7050 0.6050 0.8050 0.6050
                 0.8050 1.3700 1.2450 1.3700 1.2450 1.8200 1.8150 1.8200 1.8150 0.6200 1.9350 0.6200 ;
    END
END TLATNTSCAX16

MACRO TLATNTSCAX12
    CLASS CORE ;
    FOREIGN TLATNTSCAX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 0.8200 0.5650 1.0900 ;
        RECT  0.3050 0.7800 0.5450 1.0900 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 0.7600 1.0900 1.2050 ;
        RECT  0.9250 0.7800 1.0450 1.2500 ;
        END
    END SE
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 0.7600 1.3850 1.2500 ;
        RECT  1.2300 0.7600 1.3850 1.2200 ;
        END
    END CK
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.9250 1.3100 11.0450 2.2100 ;
        RECT  10.0850 1.0400 11.0450 1.1600 ;
        RECT  10.9250 0.4050 11.0450 1.1600 ;
        RECT  10.7450 1.3100 11.0450 1.4300 ;
        RECT  7.5850 1.1900 10.8650 1.3100 ;
        RECT  10.0850 1.0400 10.8650 1.3100 ;
        RECT  10.0850 0.4050 10.2050 2.2100 ;
        RECT  9.2450 0.4050 9.3650 2.2100 ;
        RECT  8.4050 1.0400 9.3650 1.3100 ;
        RECT  8.4050 0.4050 8.5250 2.2100 ;
        RECT  7.5850 1.1750 7.7600 1.4350 ;
        RECT  7.5850 0.8000 7.7050 1.4500 ;
        RECT  7.5650 1.3300 7.6850 2.2100 ;
        RECT  7.5650 0.4000 7.6850 0.9200 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  11.3450 -0.1800 11.4650 0.9200 ;
        RECT  10.5050 -0.1800 10.6250 0.9200 ;
        RECT  9.6650 -0.1800 9.7850 0.9200 ;
        RECT  8.8250 -0.1800 8.9450 0.9200 ;
        RECT  7.9850 -0.1800 8.1050 0.9200 ;
        RECT  7.1450 -0.1800 7.2650 0.6400 ;
        RECT  6.0450 0.4700 6.2850 0.5900 ;
        RECT  6.0450 -0.1800 6.1650 0.5900 ;
        RECT  4.7650 -0.1800 4.8850 0.5800 ;
        RECT  2.9350 0.6900 3.1750 0.8100 ;
        RECT  2.9350 -0.1800 3.0550 0.8100 ;
        RECT  1.0650 -0.1800 1.1850 0.6400 ;
        RECT  0.2250 -0.1800 0.3450 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  11.3450 1.4300 11.4650 2.7900 ;
        RECT  10.5050 1.4300 10.6250 2.7900 ;
        RECT  9.6650 1.4300 9.7850 2.7900 ;
        RECT  8.8250 1.4300 8.9450 2.7900 ;
        RECT  7.9850 1.4300 8.1050 2.7900 ;
        RECT  7.0850 1.7200 7.3250 2.1500 ;
        RECT  7.0850 1.7200 7.2050 2.7900 ;
        RECT  6.3050 1.7200 6.4250 2.7900 ;
        RECT  5.4650 1.7200 5.5850 2.7900 ;
        RECT  4.6250 1.4400 4.7450 2.7900 ;
        RECT  3.2950 2.1300 3.4150 2.7900 ;
        RECT  3.1750 2.1300 3.4150 2.2500 ;
        RECT  1.0050 1.6100 1.1250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.4650 1.2100 7.0850 1.2100 7.0850 1.6000 6.8450 1.6000 6.8450 2.2100 6.7250 2.2100
                 6.7250 1.6000 6.0050 1.6000 6.0050 2.2100 5.8850 2.2100 5.8850 1.6000 5.1650 1.6000
                 5.1650 2.0900 5.0450 2.0900 5.0450 1.4800 6.9650 1.4800 6.9650 0.8800 6.7450 0.8800
                 6.7450 0.8300 5.5250 0.8300 5.5250 0.7800 5.4050 0.7800 5.4050 0.6600 5.6450 0.6600
                 5.6450 0.7100 6.7450 0.7100 6.7450 0.6000 6.8650 0.6000 6.8650 0.7600 7.0850 0.7600
                 7.0850 1.0900 7.4650 1.0900 ;
        POLYGON  6.8450 1.1200 5.1650 1.1200 5.1650 0.8200 4.5250 0.8200 4.5250 0.4800 3.7750 0.4800
                 3.7750 0.7600 3.7350 0.7600 3.7350 1.2900 3.0750 1.2900 3.0750 1.6500 3.8950 1.6500
                 3.8950 1.8900 4.0150 1.8900 4.0150 2.0100 3.7750 2.0100 3.7750 1.7700 2.9550 1.7700
                 2.9550 1.3700 2.8350 1.3700 2.8350 1.1700 3.6150 1.1700 3.6150 0.6400 3.6550 0.6400
                 3.6550 0.3600 4.6450 0.3600 4.6450 0.7000 5.2850 0.7000 5.2850 1.0000 6.8450 1.0000 ;
        POLYGON  6.2250 1.3600 4.9250 1.3600 4.9250 1.0600 4.2650 1.0600 4.2650 1.6800 4.1450 1.6800
                 4.1450 1.5300 3.1950 1.5300 3.1950 1.4100 4.1450 1.4100 4.1450 0.7200 4.2850 0.7200
                 4.2850 0.6000 4.4050 0.6000 4.4050 0.9400 5.0450 0.9400 5.0450 1.2400 6.2250 1.2400 ;
        POLYGON  4.6250 1.3000 4.5050 1.3000 4.5050 1.9200 4.4500 1.9200 4.4500 2.2500 3.5350 2.2500
                 3.5350 2.0100 2.6550 2.0100 2.6550 2.1100 2.5350 2.1100 2.5350 1.9900 2.3550 1.9900
                 2.3550 0.8200 2.2350 0.8200 2.2350 0.7000 2.4750 0.7000 2.4750 1.8700 2.6550 1.8700
                 2.6550 1.8900 3.6550 1.8900 3.6550 2.1300 4.3300 2.1300 4.3300 1.8000 4.3850 1.8000
                 4.3850 1.1800 4.6250 1.1800 ;
        POLYGON  3.5350 0.4800 3.4150 0.4800 3.4150 1.0500 2.7150 1.0500 2.7150 1.5100 2.7950 1.5100
                 2.7950 1.7500 2.6750 1.7500 2.6750 1.6300 2.5950 1.6300 2.5950 0.5800 2.3300 0.5800
                 2.3300 0.5200 1.6250 0.5200 1.6250 1.4900 1.6050 1.4900 1.6050 1.7300 1.4850 1.7300
                 1.4850 1.3700 1.5050 1.3700 1.5050 0.6400 1.4850 0.6400 1.4850 0.4000 2.0950 0.4000
                 2.0950 0.3800 2.3350 0.3800 2.3350 0.4000 2.4500 0.4000 2.4500 0.4600 2.8150 0.4600
                 2.8150 0.9300 3.2950 0.9300 3.2950 0.3600 3.5350 0.3600 ;
        POLYGON  2.2350 2.0700 2.1150 2.0700 2.1150 1.9700 1.2450 1.9700 1.2450 1.4900 0.4850 1.4900
                 0.4850 1.7300 0.3650 1.7300 0.3650 1.3700 0.6850 1.3700 0.6850 0.6600 0.6450 0.6600
                 0.6450 0.4000 0.7650 0.4000 0.7650 0.5400 0.8050 0.5400 0.8050 1.3700 1.3650 1.3700
                 1.3650 1.8500 1.9350 1.8500 1.9350 0.8200 1.8150 0.8200 1.8150 0.7000 2.0550 0.7000
                 2.0550 1.8300 2.2350 1.8300 ;
    END
END TLATNTSCAX12

MACRO TLATNSRXL
    CLASS CORE ;
    FOREIGN TLATNSRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9450 1.2500 2.0650 1.4900 ;
        RECT  1.7550 1.5200 2.0150 1.6700 ;
        RECT  1.8950 1.3700 2.0150 1.6700 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9800 1.1200 5.1750 1.4950 ;
        RECT  4.9800 1.1200 5.1200 1.5000 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6700 1.2550 6.9100 1.3750 ;
        RECT  6.1900 1.1750 6.7900 1.2950 ;
        RECT  6.1900 0.8850 6.4750 1.2950 ;
        RECT  6.3550 0.3750 6.4750 1.2950 ;
        RECT  5.4250 0.3750 6.4750 0.4950 ;
        RECT  6.1600 0.8850 6.4750 1.1450 ;
        RECT  4.7750 0.6400 5.5450 0.7600 ;
        RECT  5.4250 0.3750 5.5450 0.7600 ;
        RECT  4.7750 0.3600 4.8950 0.7600 ;
        RECT  3.0650 0.3600 4.8950 0.4800 ;
        END
    END RN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0300 1.1750 7.3350 1.4150 ;
        RECT  7.0300 1.1750 7.1800 1.4350 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 1.5850 1.4850 1.8300 ;
        RECT  1.3650 0.6500 1.4850 0.8900 ;
        RECT  1.2300 1.4650 1.4450 1.7250 ;
        RECT  1.3250 0.7700 1.4450 1.7250 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  7.1550 -0.1800 7.2750 0.7950 ;
        RECT  5.1850 -0.1800 5.3050 0.5200 ;
        RECT  2.8250 0.6800 3.1650 0.8000 ;
        RECT  2.8250 -0.1800 2.9450 0.8000 ;
        RECT  1.7850 -0.1800 1.9050 0.8900 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  7.0300 1.6550 7.1500 2.7900 ;
        RECT  6.1900 1.6550 6.3100 2.7900 ;
        RECT  5.0650 1.6200 5.1850 2.7900 ;
        RECT  3.5250 1.8900 3.6450 2.7900 ;
        RECT  2.6850 2.2300 2.8050 2.7900 ;
        RECT  1.8450 2.2300 1.9650 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.6950 0.9350 7.5750 0.9350 7.5750 1.6550 7.5700 1.6550 7.5700 1.7750 7.4500 1.7750
                 7.4500 1.5350 7.4550 1.5350 7.4550 1.0550 6.5950 1.0550 6.5950 0.9350 7.4550 0.9350
                 7.4550 0.8150 7.5750 0.8150 7.5750 0.5550 7.6950 0.5550 ;
        POLYGON  6.7300 1.7750 6.6100 1.7750 6.6100 1.6550 6.4300 1.6550 6.4300 1.5350 5.9200 1.5350
                 5.9200 1.2400 5.5450 1.2400 5.5450 1.1200 5.9200 1.1200 5.9200 0.6150 6.2350 0.6150
                 6.2350 0.7350 6.0400 0.7350 6.0400 1.4150 6.5500 1.4150 6.5500 1.5350 6.7300 1.5350 ;
        POLYGON  5.7850 1.0000 5.4250 1.0000 5.4250 1.5000 5.6050 1.5000 5.6050 1.7400 5.4850 1.7400
                 5.4850 1.6200 5.3050 1.6200 5.3050 1.0000 4.8450 1.0000 4.8450 1.1200 4.1850 1.1200
                 4.1850 1.2000 3.9450 1.2000 3.9450 1.0800 4.0650 1.0800 4.0650 1.0000 4.7250 1.0000
                 4.7250 0.8800 5.6650 0.8800 5.6650 0.6200 5.7850 0.6200 ;
        POLYGON  4.6050 0.8800 3.8250 0.8800 3.8250 1.3200 4.4450 1.3200 4.4450 1.7400 4.3250 1.7400
                 4.3250 1.4400 2.4250 1.4400 2.4250 1.3200 3.7050 1.3200 3.7050 0.7600 4.4850 0.7600
                 4.4850 0.6200 4.6050 0.6200 ;
        POLYGON  4.0850 1.6800 3.9650 1.6800 3.9650 1.7700 2.9850 1.7700 2.9850 1.6500 3.8450 1.6500
                 3.8450 1.5600 4.0850 1.5600 ;
        POLYGON  3.5850 1.2000 3.4650 1.2000 3.4650 1.1300 2.3050 1.1300 2.3050 1.5900 2.3250 1.5900
                 2.3250 1.8300 2.2050 1.8300 2.2050 1.7100 2.1850 1.7100 2.1850 1.1300 1.8050 1.1300
                 1.8050 1.1700 1.5650 1.1700 1.5650 1.0100 2.4250 1.0100 2.4250 0.6500 2.5450 0.6500
                 2.5450 1.0100 3.4650 1.0100 3.4650 0.9600 3.5850 0.9600 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END TLATNSRXL

MACRO TLATNSRX4
    CLASS CORE ;
    FOREIGN TLATNSRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1400 0.5200 1.5900 ;
        END
    END GN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1900 0.4000 4.7550 0.5200 ;
        RECT  2.1300 0.5000 3.3100 0.6200 ;
        RECT  2.1300 0.3600 2.2500 0.6200 ;
        RECT  1.3550 0.3600 2.2500 0.4800 ;
        RECT  0.6550 1.1600 1.4750 1.2800 ;
        RECT  1.3550 0.3600 1.4750 1.2800 ;
        RECT  1.1750 1.1600 1.4350 1.3800 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.4650 2.6700 1.5850 ;
        RECT  2.5500 1.3350 2.6700 1.5850 ;
        RECT  2.3900 1.4650 2.5400 1.7300 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8150 1.1500 6.3950 1.2700 ;
        RECT  5.8150 1.1500 6.0750 1.3800 ;
        RECT  5.2550 1.3600 5.9350 1.4800 ;
        RECT  5.2550 1.1700 5.3750 1.4800 ;
        RECT  5.0950 1.1700 5.3750 1.2900 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8550 1.3100 7.9750 2.0800 ;
        RECT  7.6750 1.3100 7.9750 1.4300 ;
        RECT  7.0350 0.8500 7.8150 0.9700 ;
        RECT  7.6950 0.6800 7.8150 0.9700 ;
        RECT  7.0300 1.1900 7.7950 1.3100 ;
        RECT  7.0300 1.1750 7.1800 1.4350 ;
        RECT  7.0350 0.8000 7.1550 1.4350 ;
        RECT  7.0150 1.3100 7.1350 2.0800 ;
        RECT  6.8550 0.8000 7.1550 0.9200 ;
        RECT  6.8550 0.6800 6.9750 0.9200 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.2150 1.3100 11.3350 2.0800 ;
        RECT  11.0350 1.3100 11.3350 1.4300 ;
        RECT  10.3950 0.8500 11.1750 0.9700 ;
        RECT  11.0550 0.6800 11.1750 0.9700 ;
        RECT  10.3950 1.1900 11.1550 1.3100 ;
        RECT  10.3950 0.8500 10.7150 1.3100 ;
        RECT  10.3750 1.3100 10.5150 1.4300 ;
        RECT  10.3750 1.3100 10.4950 2.0800 ;
        RECT  10.2150 0.8000 10.5150 0.9200 ;
        RECT  10.2150 0.6800 10.3350 0.9200 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  11.4750 -0.1800 11.5950 0.7300 ;
        RECT  10.6350 -0.1800 10.7550 0.7300 ;
        RECT  9.7950 -0.1800 9.9150 0.7300 ;
        RECT  8.9550 -0.1800 9.0750 0.7300 ;
        RECT  8.1150 -0.1800 8.2350 0.7300 ;
        RECT  7.2750 -0.1800 7.3950 0.7300 ;
        RECT  6.4350 -0.1800 6.5550 0.7300 ;
        RECT  5.0150 -0.1800 5.1350 0.8000 ;
        RECT  2.9150 -0.1800 3.0350 0.3800 ;
        RECT  2.5250 -0.1800 2.6450 0.3800 ;
        RECT  0.5550 -0.1800 0.6750 0.7800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  11.6350 1.4300 11.7550 2.7900 ;
        RECT  10.7950 1.4300 10.9150 2.7900 ;
        RECT  9.9550 1.4300 10.0750 2.7900 ;
        RECT  9.1150 1.4300 9.2350 2.7900 ;
        RECT  8.2750 1.4300 8.3950 2.7900 ;
        RECT  7.4350 1.4300 7.5550 2.7900 ;
        RECT  6.5950 1.8400 6.7150 2.7900 ;
        RECT  5.7550 2.2300 5.8750 2.7900 ;
        RECT  4.9150 2.2300 5.0350 2.7900 ;
        RECT  3.9550 2.0000 4.0750 2.7900 ;
        RECT  2.2700 2.2200 2.5100 2.7900 ;
        RECT  1.4000 2.2200 1.6400 2.7900 ;
        RECT  0.5000 2.2300 0.6200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.2750 1.1800 9.4750 1.1800 9.4750 1.3100 9.6550 1.3100 9.6550 2.0800 9.5350 2.0800
                 9.5350 1.4300 9.3550 1.4300 9.3550 1.3100 8.8150 1.3100 8.8150 2.0800 8.6950 2.0800
                 8.6950 0.9200 8.5350 0.9200 8.5350 0.6800 8.6550 0.6800 8.6550 0.8000 8.8150 0.8000
                 8.8150 1.0600 9.3750 1.0600 9.3750 0.6800 9.4950 0.6800 9.4950 1.0600 10.2750 1.0600 ;
        POLYGON  6.7350 1.2400 6.6350 1.2400 6.6350 1.7200 6.2350 1.7200 6.2350 1.9500 6.1150 1.9500
                 6.1150 1.7200 5.3950 1.7200 5.3950 1.9500 5.2750 1.9500 5.2750 1.7200 4.8550 1.7200
                 4.8550 1.4500 4.2950 1.4500 4.2950 1.3300 4.9750 1.3300 4.9750 1.6000 6.5150 1.6000
                 6.5150 1.0300 5.7350 1.0300 5.7350 0.6600 5.8550 0.6600 5.8550 0.9100 6.7350 0.9100 ;
        POLYGON  5.6150 1.2400 5.4950 1.2400 5.4950 1.0400 4.1750 1.0400 4.1750 1.6400 3.2300 1.6400
                 3.2300 1.8200 3.1500 1.8200 3.1500 1.9400 3.0300 1.9400 3.0300 1.7000 3.1100 1.7000
                 3.1100 1.5200 4.0550 1.5200 4.0550 1.0400 3.6950 1.0400 3.6950 0.9200 3.6150 0.9200
                 3.6150 0.6600 3.7350 0.6600 3.7350 0.8000 3.8150 0.8000 3.8150 0.9200 5.6150 0.9200 ;
        RECT  3.3900 1.7600 4.6150 1.8800 ;
        POLYGON  3.9350 1.2800 3.8150 1.2800 3.8150 1.4000 2.9900 1.4000 2.9900 1.5800 2.9100 1.5800
                 2.9100 1.9700 2.2700 1.9700 2.2700 2.1000 1.5500 2.1000 1.5500 1.6200 1.1000 1.6200
                 1.1000 1.8300 0.9800 1.8300 0.9800 1.5000 1.5950 1.5000 1.5950 0.6000 1.8350 0.6000
                 1.8350 0.7200 1.7150 0.7200 1.7150 1.6200 1.6700 1.6200 1.6700 1.9800 2.1500 1.9800
                 2.1500 1.2250 2.3900 1.2250 2.3900 1.3450 2.2700 1.3450 2.2700 1.8500 2.7900 1.8500
                 2.7900 1.2800 3.6950 1.2800 3.6950 1.1600 3.9350 1.1600 ;
        POLYGON  3.5750 1.1600 3.3350 1.1600 3.3350 1.1050 2.0300 1.1050 2.0300 1.8600 1.7900 1.8600
                 1.7900 1.7400 1.9100 1.7400 1.9100 0.8400 1.9850 0.8400 1.9850 0.7400 2.2250 0.7400
                 2.2250 0.9850 3.4550 0.9850 3.4550 1.0400 3.5750 1.0400 ;
        POLYGON  1.2350 1.0400 0.9950 1.0400 0.9950 1.0200 0.2400 1.0200 0.2400 1.7100 0.2550 1.7100
                 0.2550 1.9500 0.1350 1.9500 0.1350 1.8300 0.1200 1.8300 0.1200 0.7800 0.1350 0.7800
                 0.1350 0.5400 0.2550 0.5400 0.2550 0.9000 1.2350 0.9000 ;
    END
END TLATNSRX4

MACRO TLATNSRX2
    CLASS CORE ;
    FOREIGN TLATNSRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6150 1.1600 0.8350 1.5100 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.3300 3.1200 1.7250 ;
        RECT  2.8800 1.3300 3.1200 1.4500 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6900 1.0900 4.8600 1.5000 ;
        RECT  4.6900 1.0900 4.8100 1.5150 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6700 1.0000 7.8100 1.2700 ;
        RECT  7.6100 0.8600 7.7800 1.1450 ;
        END
    END GN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3300 0.6800 5.4500 1.0250 ;
        RECT  5.2700 1.3800 5.3900 1.6700 ;
        RECT  5.3200 0.8850 5.4400 1.5000 ;
        RECT  5.2900 0.8850 5.4400 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.1900 1.1450 7.3100 1.6700 ;
        RECT  7.0600 1.1450 7.3100 1.2650 ;
        RECT  7.0300 0.8850 7.1800 1.1450 ;
        RECT  7.0100 0.6800 7.1300 1.0250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.4300 -0.1800 7.5500 0.7300 ;
        RECT  6.5900 -0.1800 6.7100 0.7300 ;
        RECT  5.7500 -0.1800 5.8700 0.7300 ;
        RECT  4.9100 -0.1800 5.0300 0.7300 ;
        RECT  2.7150 0.6100 2.9550 0.7300 ;
        RECT  2.7150 -0.1800 2.8350 0.7300 ;
        RECT  0.4950 0.6800 0.7350 0.8000 ;
        RECT  0.4950 -0.1800 0.6150 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.6700 2.0300 7.7900 2.7900 ;
        RECT  6.6500 2.0300 6.8900 2.1500 ;
        RECT  6.6500 2.0300 6.7700 2.7900 ;
        RECT  5.6900 2.0300 5.9300 2.1500 ;
        RECT  5.6900 2.0300 5.8100 2.7900 ;
        RECT  4.7900 2.2300 4.9100 2.7900 ;
        RECT  4.2900 2.2300 4.4100 2.7900 ;
        RECT  3.1500 2.2300 3.2700 2.7900 ;
        RECT  2.2450 2.2900 2.4850 2.7900 ;
        RECT  0.6150 1.8700 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2700 1.7900 7.8800 1.7900 7.8800 1.9100 5.4950 1.9100 5.4950 2.1100 4.1700 2.1100
                 4.1700 2.2500 3.6100 2.2500 3.6100 2.1300 4.0500 2.1300 4.0500 1.9900 5.3750 1.9900
                 5.3750 1.7900 7.7600 1.7900 7.7600 1.6700 8.1500 1.6700 8.1500 1.5500 7.9300 1.5500
                 7.9300 0.6800 8.0500 0.6800 8.0500 1.4300 8.2700 1.4300 ;
        POLYGON  6.9100 1.2900 6.3500 1.2900 6.3500 1.6700 6.2300 1.6700 6.2300 0.9200 6.1700 0.9200
                 6.1700 0.6800 6.2900 0.6800 6.2900 0.8000 6.3500 0.8000 6.3500 1.1700 6.9100 1.1700 ;
        POLYGON  5.1700 1.2600 5.0500 1.2600 5.0500 0.9700 4.5500 0.9700 4.5500 1.8700 4.4300 1.8700
                 4.4300 0.9700 4.2100 0.9700 4.2100 0.5800 3.9450 0.5800 3.9450 0.5000 3.2700 0.5000
                 3.2700 0.9700 2.2750 0.9700 2.2750 0.4800 2.1550 0.4800 2.1550 0.3600 2.3950 0.3600
                 2.3950 0.8500 3.1500 0.8500 3.1500 0.3800 4.0650 0.3800 4.0650 0.4600 4.3300 0.4600
                 4.3300 0.8500 5.1700 0.8500 ;
        POLYGON  4.2700 1.8700 3.9300 1.8700 3.9300 2.0100 3.2050 2.0100 3.2050 2.1100 2.9400 2.1100
                 2.9400 2.1700 1.4950 2.1700 1.4950 1.7500 1.6150 1.7500 1.6150 1.5700 1.6550 1.5700
                 1.6550 0.6200 1.7750 0.6200 1.7750 1.6900 1.7350 1.6900 1.7350 1.8700 1.6150 1.8700
                 1.6150 2.0500 2.8200 2.0500 2.8200 1.9900 3.0850 1.9900 3.0850 1.8900 3.8100 1.8900
                 3.8100 1.7500 4.1500 1.7500 4.1500 1.1100 4.2700 1.1100 ;
        POLYGON  3.6900 1.7700 3.4500 1.7700 3.4500 1.2100 1.9150 1.2100 1.9150 0.5000 1.5350 0.5000
                 1.5350 1.4500 1.4150 1.4500 1.4150 1.0400 0.4950 1.0400 0.4950 1.2200 0.3550 1.2200
                 0.3550 0.9800 0.3750 0.9800 0.3750 0.9200 1.4150 0.9200 1.4150 0.3800 2.0350 0.3800
                 2.0350 1.0200 2.1550 1.0200 2.1550 1.0900 3.4750 1.0900 3.4750 0.6200 3.5950 0.6200
                 3.5950 1.2100 3.5700 1.2100 3.5700 1.6500 3.6900 1.6500 ;
        POLYGON  2.8500 1.8700 2.0950 1.8700 2.0950 1.9300 1.8550 1.9300 1.8550 1.8100 1.9750 1.8100
                 1.9750 1.7500 2.8500 1.7500 ;
        POLYGON  1.2350 1.2800 1.0750 1.2800 1.0750 1.7500 0.3150 1.7500 0.3150 1.9900 0.1950 1.9900
                 0.1950 1.8700 0.1150 1.8700 0.1150 0.7400 0.1350 0.7400 0.1350 0.6200 0.2550 0.6200
                 0.2550 0.8600 0.2350 0.8600 0.2350 1.6300 0.9550 1.6300 0.9550 1.1600 1.2350 1.1600 ;
    END
END TLATNSRX2

MACRO TLATNSRX1
    CLASS CORE ;
    FOREIGN TLATNSRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8450 1.3000 2.1650 1.4200 ;
        RECT  1.8100 1.4650 1.9650 1.7250 ;
        RECT  1.8450 1.3000 1.9650 1.7250 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 1.1750 5.1500 1.5100 ;
        RECT  4.9150 1.2400 5.0350 1.5700 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6700 1.4000 6.9100 1.5200 ;
        RECT  6.2450 1.3600 6.7900 1.4800 ;
        RECT  6.1050 1.2300 6.3750 1.3800 ;
        RECT  6.2550 0.4800 6.3750 1.4800 ;
        RECT  5.2650 0.4800 6.3750 0.6000 ;
        RECT  4.7250 0.5000 5.3850 0.6200 ;
        RECT  3.0150 0.4000 4.8450 0.5200 ;
        END
    END RN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.1550 1.2800 7.2750 1.5650 ;
        RECT  7.0300 1.4300 7.1800 1.7250 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 2.2100 ;
        RECT  1.2300 1.1750 1.4850 1.4350 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  6.9950 -0.1800 7.1150 0.9200 ;
        RECT  5.0250 -0.1800 5.1450 0.3800 ;
        RECT  2.7750 0.7200 3.1150 0.8400 ;
        RECT  2.7750 -0.1800 2.8950 0.8400 ;
        RECT  1.7850 -0.1800 1.9050 0.7300 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  6.9950 1.8450 7.1150 2.7900 ;
        RECT  6.1550 1.8450 6.2750 2.7900 ;
        RECT  5.0750 1.7000 5.1950 2.7900 ;
        RECT  3.5850 2.0700 3.7050 2.7900 ;
        RECT  2.7450 2.2300 2.8650 2.7900 ;
        RECT  1.7850 1.8450 1.9050 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.5350 1.9650 7.4150 1.9650 7.4150 1.1600 6.6150 1.1600 6.6150 1.2400 6.4950 1.2400
                 6.4950 1.0000 6.6150 1.0000 6.6150 1.0400 7.4150 1.0400 7.4150 0.6800 7.5350 0.6800 ;
        POLYGON  6.6950 1.9650 6.5750 1.9650 6.5750 1.8450 6.4300 1.8450 6.4300 1.7250 5.8650 1.7250
                 5.8650 1.3400 5.5100 1.3400 5.5100 1.2200 5.8650 1.2200 5.8650 0.7400 6.1350 0.7400
                 6.1350 0.8600 5.9850 0.8600 5.9850 1.6050 6.5500 1.6050 6.5500 1.7250 6.6950 1.7250 ;
        POLYGON  5.7450 0.8400 5.6250 0.8400 5.6250 1.0550 5.3900 1.0550 5.3900 1.4600 5.6150 1.4600
                 5.6150 1.8200 5.4950 1.8200 5.4950 1.5800 5.2700 1.5800 5.2700 1.0550 4.7950 1.0550
                 4.7950 1.3800 3.9750 1.3800 3.9750 1.2600 4.5950 1.2600 4.5950 1.0200 4.6750 1.0200
                 4.6750 0.9350 5.5050 0.9350 5.5050 0.7200 5.7450 0.7200 ;
        POLYGON  4.5550 0.9000 4.4750 0.9000 4.4750 1.1400 3.8550 1.1400 3.8550 1.5000 4.4350 1.5000
                 4.4350 1.8200 4.3150 1.8200 4.3150 1.6200 3.7350 1.6200 3.7350 1.5100 2.5450 1.5100
                 2.5450 1.2700 2.6650 1.2700 2.6650 1.3900 3.7350 1.3900 3.7350 1.0200 4.3550 1.0200
                 4.3550 0.7800 4.4350 0.7800 4.4350 0.6600 4.5550 0.6600 ;
        RECT  3.0450 1.7400 4.0750 1.8600 ;
        POLYGON  3.6150 1.1600 3.3750 1.1600 3.3750 1.1500 2.4050 1.1500 2.4050 1.6600 2.3850 1.6600
                 2.3850 1.8300 2.2650 1.8300 2.2650 1.5400 2.2850 1.5400 2.2850 1.1500 1.7250 1.1500
                 1.7250 1.2700 1.6050 1.2700 1.6050 1.0300 2.4850 1.0300 2.4850 0.6800 2.6050 0.6800
                 2.6050 1.0300 3.6150 1.0300 ;
        POLYGON  1.0950 1.9900 0.9750 1.9900 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END TLATNSRX1

MACRO TLATNCAX8
    CLASS CORE ;
    FOREIGN TLATNCAX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.4650 0.5650 1.6700 ;
        RECT  0.4450 1.2600 0.5650 1.6700 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.5150 1.1450 1.7200 ;
        RECT  0.9150 1.3600 1.0350 1.7200 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1550 1.1000 8.2750 2.0800 ;
        RECT  8.1350 0.6450 8.2550 1.2200 ;
        RECT  5.6100 1.1000 8.2750 1.2200 ;
        RECT  6.5150 0.7650 8.2550 0.8850 ;
        RECT  7.2350 0.7150 7.4750 0.8850 ;
        RECT  7.3150 1.1000 7.4350 2.0800 ;
        RECT  6.3950 0.7150 6.6350 0.8350 ;
        RECT  6.4750 1.1000 6.5950 2.0850 ;
        RECT  5.6350 1.1000 5.7550 2.0850 ;
        RECT  5.5550 0.8850 5.7300 1.1000 ;
        RECT  5.5550 0.6550 5.6750 1.1000 ;
        RECT  5.6100 1.1000 5.7550 1.3400 ;
        RECT  5.5800 1.1000 8.2750 1.1450 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.7150 -0.1800 7.8350 0.6450 ;
        RECT  6.8750 -0.1800 6.9950 0.6450 ;
        RECT  5.9750 -0.1800 6.0950 0.6400 ;
        RECT  5.1350 -0.1800 5.2550 0.6400 ;
        RECT  3.7350 0.4500 3.9750 0.5700 ;
        RECT  3.8550 -0.1800 3.9750 0.5700 ;
        RECT  2.2750 -0.1800 2.3950 0.3800 ;
        RECT  0.5550 -0.1800 0.6750 0.9000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.7350 1.3400 7.8550 2.7900 ;
        RECT  6.8950 1.3400 7.0150 2.7900 ;
        RECT  6.0550 1.3400 6.1750 2.7900 ;
        RECT  5.2150 1.7700 5.3350 2.7900 ;
        RECT  4.3750 1.7700 4.4950 2.7900 ;
        RECT  3.4750 2.2300 3.5950 2.7900 ;
        RECT  2.0750 2.2600 2.3150 2.7900 ;
        RECT  0.7550 1.8400 0.8750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.4350 1.2150 5.3350 1.2150 5.3350 1.6500 4.9150 1.6500 4.9150 2.0800 4.7950 2.0800
                 4.7950 1.6500 4.0750 1.6500 4.0750 2.0800 3.9550 2.0800 3.9550 1.5300 5.2150 1.5300
                 5.2150 0.9700 4.5750 0.9700 4.5750 0.8100 4.4950 0.8100 4.4950 0.5700 4.6150 0.5700
                 4.6150 0.6900 4.6950 0.6900 4.6950 0.8500 5.4350 0.8500 ;
        POLYGON  5.0950 1.4100 3.8750 1.4100 3.8750 1.0500 3.2550 1.0500 3.2550 1.4300 3.1250 1.4300
                 3.1250 1.8700 3.0050 1.8700 3.0050 1.4300 2.0750 1.4300 2.0750 1.3100 3.1350 1.3100
                 3.1350 0.6500 3.3750 0.6500 3.3750 0.7700 3.2550 0.7700 3.2550 0.9300 3.9950 0.9300
                 3.9950 1.2900 4.9750 1.2900 4.9750 1.0900 5.0950 1.0900 ;
        POLYGON  4.4550 1.1700 4.3350 1.1700 4.3350 1.0500 4.2550 1.0500 4.2550 0.8100 3.4950 0.8100
                 3.4950 0.5300 3.0150 0.5300 3.0150 0.7400 2.8750 0.7400 2.8750 1.1800 1.9550 1.1800
                 1.9550 1.7400 2.6750 1.7400 2.6750 1.7800 2.7950 1.7800 2.7950 1.9000 2.5550 1.9000
                 2.5550 1.8600 1.8350 1.8600 1.8350 1.1800 1.7550 1.1800 1.7550 1.0600 2.7550 1.0600
                 2.7550 0.6200 2.8950 0.6200 2.8950 0.4100 3.6150 0.4100 3.6150 0.6900 4.3750 0.6900
                 4.3750 0.9300 4.4550 0.9300 ;
        POLYGON  3.6150 1.2900 3.4950 1.2900 3.4950 2.1100 3.1450 2.1100 3.1450 2.1400 2.2300 2.1400
                 2.2300 2.1000 1.4350 2.1000 1.4350 1.8600 1.2750 1.8600 1.2750 0.6600 1.3950 0.6600
                 1.3950 1.7400 1.5550 1.7400 1.5550 1.9800 2.3500 1.9800 2.3500 2.0200 3.0250 2.0200
                 3.0250 1.9900 3.3750 1.9900 3.3750 1.1700 3.6150 1.1700 ;
        POLYGON  2.7750 0.5000 2.6350 0.5000 2.6350 0.6200 2.0350 0.6200 2.0350 0.5400 1.6350 0.5400
                 1.6350 1.3800 1.7150 1.3800 1.7150 1.6200 1.5150 1.6200 1.5150 0.5400 1.1550 0.5400
                 1.1550 1.2400 1.0350 1.2400 1.0350 1.1400 0.1850 1.1400 0.1850 1.7900 0.4550 1.7900
                 0.4550 2.0300 0.3350 2.0300 0.3350 1.9100 0.0650 1.9100 0.0650 0.9000 0.1350 0.9000
                 0.1350 0.6600 0.2550 0.6600 0.2550 1.0200 1.0350 1.0200 1.0350 0.4200 2.1550 0.4200
                 2.1550 0.5000 2.5150 0.5000 2.5150 0.3800 2.7750 0.3800 ;
    END
END TLATNCAX8

MACRO TLATNCAX6
    CLASS CORE ;
    FOREIGN TLATNCAX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4450 1.1400 0.5650 1.5200 ;
        RECT  0.3050 1.1650 0.5650 1.3800 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.4650 1.1450 1.6700 ;
        RECT  0.9350 1.3600 1.0550 1.7100 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2850 1.3400 7.4050 2.1200 ;
        RECT  7.2650 0.4050 7.3850 1.0400 ;
        RECT  7.1050 1.3400 7.4050 1.4600 ;
        RECT  7.0850 0.9200 7.3850 1.0400 ;
        RECT  7.1050 0.9200 7.2250 1.4600 ;
        RECT  5.6050 1.0400 7.2250 1.1600 ;
        RECT  6.4450 1.0400 6.5650 2.1200 ;
        RECT  6.4250 0.4050 6.5450 1.1600 ;
        RECT  5.5250 0.8850 5.7300 1.0400 ;
        RECT  5.6050 0.8850 5.7250 2.1200 ;
        RECT  5.5250 0.4000 5.6450 1.0400 ;
        RECT  5.5800 1.0400 7.2250 1.1450 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.8450 -0.1800 6.9650 0.9200 ;
        RECT  6.0050 -0.1800 6.1250 0.9200 ;
        RECT  5.1050 -0.1800 5.2250 0.7300 ;
        RECT  3.7050 0.4500 3.9450 0.5700 ;
        RECT  3.8250 -0.1800 3.9450 0.5700 ;
        RECT  2.2450 -0.1800 2.3650 0.3800 ;
        RECT  0.6150 -0.1800 0.7350 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.8650 1.3400 6.9850 2.7900 ;
        RECT  6.0250 1.3400 6.1450 2.7900 ;
        RECT  5.1850 1.7700 5.3050 2.7900 ;
        RECT  4.3450 1.7700 4.4650 2.7900 ;
        RECT  3.4450 2.2300 3.5650 2.7900 ;
        RECT  2.0550 2.2500 2.2950 2.7900 ;
        RECT  0.7550 1.8300 0.8750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.4050 1.2400 5.3050 1.2400 5.3050 1.6500 4.8850 1.6500 4.8850 2.0800 4.7650 2.0800
                 4.7650 1.6500 4.0450 1.6500 4.0450 2.0800 3.9250 2.0800 3.9250 1.5300 5.1850 1.5300
                 5.1850 0.9700 4.5450 0.9700 4.5450 0.8100 4.4650 0.8100 4.4650 0.5700 4.5850 0.5700
                 4.5850 0.6900 4.6650 0.6900 4.6650 0.8500 5.4050 0.8500 ;
        POLYGON  5.0650 1.4100 3.7650 1.4100 3.7650 1.0500 3.2250 1.0500 3.2250 1.3700 3.1050 1.3700
                 3.1050 1.8700 2.9850 1.8700 2.9850 1.3700 2.0550 1.3700 2.0550 1.2500 3.1050 1.2500
                 3.1050 0.6500 3.3450 0.6500 3.3450 0.7700 3.2250 0.7700 3.2250 0.9300 3.8850 0.9300
                 3.8850 1.2900 4.9450 1.2900 4.9450 1.0900 5.0650 1.0900 ;
        POLYGON  4.4250 1.1700 4.3050 1.1700 4.3050 1.0500 4.2250 1.0500 4.2250 0.8100 3.4650 0.8100
                 3.4650 0.5300 2.9850 0.5300 2.9850 0.7800 2.8450 0.7800 2.8450 1.1300 1.9350 1.1300
                 1.9350 1.7300 2.6450 1.7300 2.6450 1.7700 2.7750 1.7700 2.7750 1.8900 2.5250 1.8900
                 2.5250 1.8500 1.8150 1.8500 1.8150 1.2500 1.7550 1.2500 1.7550 1.0100 2.7250 1.0100
                 2.7250 0.6600 2.8650 0.6600 2.8650 0.4100 3.5850 0.4100 3.5850 0.6900 4.3450 0.6900
                 4.3450 0.9300 4.4250 0.9300 ;
        POLYGON  3.5850 1.2900 3.4650 1.2900 3.4650 2.1100 3.2000 2.1100 3.2000 2.1300 2.2850 2.1300
                 2.2850 2.0900 1.4150 2.0900 1.4150 1.8500 1.2750 1.8500 1.2750 0.6600 1.3950 0.6600
                 1.3950 1.7300 1.5350 1.7300 1.5350 1.9700 2.4050 1.9700 2.4050 2.0100 3.0800 2.0100
                 3.0800 1.9900 3.3450 1.9900 3.3450 1.1700 3.5850 1.1700 ;
        POLYGON  2.7450 0.5000 2.6050 0.5000 2.6050 0.6200 2.0050 0.6200 2.0050 0.5400 1.6350 0.5400
                 1.6350 1.3700 1.6950 1.3700 1.6950 1.6100 1.5750 1.6100 1.5750 1.4900 1.5150 1.4900
                 1.5150 0.5400 1.1550 0.5400 1.1550 1.2400 1.0350 1.2400 1.0350 1.0200 0.1850 1.0200
                 0.1850 1.6400 0.4550 1.6400 0.4550 1.9500 0.3350 1.9500 0.3350 1.7600 0.0650 1.7600
                 0.0650 0.7800 0.1350 0.7800 0.1350 0.6600 0.2550 0.6600 0.2550 0.9000 1.0350 0.9000
                 1.0350 0.4200 2.1250 0.4200 2.1250 0.5000 2.4850 0.5000 2.4850 0.3800 2.7450 0.3800 ;
    END
END TLATNCAX6

MACRO TLATNCAX4
    CLASS CORE ;
    FOREIGN TLATNCAX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8850 0.8350 1.1850 ;
        RECT  0.6100 0.9550 0.7700 1.2400 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5250 1.2200 5.7850 1.4400 ;
        RECT  5.5250 1.2200 5.6450 1.5700 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0350 1.4000 2.2750 1.5800 ;
        RECT  2.0150 0.7400 2.2550 0.8600 ;
        RECT  1.2350 0.7900 2.1350 0.9100 ;
        RECT  1.2300 1.3000 2.1550 1.4200 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        RECT  1.2350 0.6700 1.3550 1.4600 ;
        RECT  1.1350 1.3400 1.2550 1.5800 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.5250 0.5000 5.7650 0.6200 ;
        RECT  5.6450 -0.1800 5.7650 0.6200 ;
        RECT  4.0050 0.6200 4.1250 0.8600 ;
        RECT  3.9650 -0.1800 4.0850 0.7400 ;
        RECT  2.4950 -0.1800 2.6150 0.7300 ;
        RECT  1.5950 0.5500 1.8350 0.6700 ;
        RECT  1.5950 -0.1800 1.7150 0.6700 ;
        RECT  0.8150 -0.1800 0.9350 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.6050 1.6900 5.7250 2.7900 ;
        RECT  4.2050 2.1000 4.4450 2.2200 ;
        RECT  4.2050 2.1000 4.3250 2.7900 ;
        RECT  3.3050 2.1200 3.4250 2.7900 ;
        RECT  2.5750 2.1200 2.6950 2.7900 ;
        RECT  1.5550 1.9400 1.7950 2.0600 ;
        RECT  1.5550 1.9400 1.6750 2.7900 ;
        RECT  0.6550 1.9400 0.7750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.2650 1.7500 5.9650 1.7500 5.9650 1.6300 6.1450 1.6300 6.1450 0.8600 5.2850 0.8600
                 5.2850 0.4800 4.2050 0.4800 4.2050 0.3600 5.4050 0.3600 5.4050 0.7400 6.0650 0.7400
                 6.0650 0.6200 6.1850 0.6200 6.1850 0.7400 6.2650 0.7400 ;
        POLYGON  6.0250 1.2200 5.9050 1.2200 5.9050 1.1000 5.4050 1.1000 5.4050 1.7100 5.1450 1.7100
                 5.1450 1.7500 4.9050 1.7500 4.9050 1.6300 5.0250 1.6300 5.0250 1.5900 5.2850 1.5900
                 5.2850 1.1000 4.7650 1.1000 4.7650 0.6200 4.8850 0.6200 4.8850 0.9800 6.0250 0.9800 ;
        POLYGON  5.1650 1.4700 5.0450 1.4700 5.0450 1.3500 3.2350 1.3500 3.2350 1.5200 2.9950 1.5200
                 2.9950 1.4000 3.1150 1.4000 3.1150 0.9200 2.9750 0.9200 2.9750 0.6800 3.0950 0.6800
                 3.0950 0.8000 3.2350 0.8000 3.2350 1.2300 4.5050 1.2300 4.5050 0.9600 4.6250 0.9600
                 4.6250 1.2300 5.1650 1.2300 ;
        POLYGON  4.9450 2.2500 4.8250 2.2500 4.8250 1.9900 4.5650 1.9900 4.5650 1.9800 3.8900 1.9800
                 3.8900 2.0000 2.4450 2.0000 2.4450 1.8200 0.1750 1.8200 0.1750 1.4600 0.3350 1.4600
                 0.3350 0.6800 0.4550 0.6800 0.4550 1.5800 0.2950 1.5800 0.2950 1.7000 2.5650 1.7000
                 2.5650 1.8800 3.7700 1.8800 3.7700 1.8600 4.6850 1.8600 4.6850 1.8700 4.9450 1.8700 ;
        POLYGON  3.9650 1.7400 3.5800 1.7400 3.5800 1.7600 2.7350 1.7600 2.7350 1.1800 1.8950 1.1800
                 1.8950 1.0600 2.7350 1.0600 2.7350 0.4400 3.4850 0.4400 3.4850 0.7300 3.3650 0.7300
                 3.3650 0.5600 2.8550 0.5600 2.8550 1.6400 3.4600 1.6400 3.4600 1.6200 3.9650 1.6200 ;
    END
END TLATNCAX4

MACRO TLATNCAX3
    CLASS CORE ;
    FOREIGN TLATNCAX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2750 1.0200 0.3950 1.2800 ;
        RECT  0.0700 1.0200 0.3950 1.1600 ;
        RECT  0.0700 0.8850 0.2200 1.1600 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3250 1.2300 1.4450 1.5800 ;
        RECT  1.1750 1.2300 1.4450 1.4350 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8250 1.3200 5.9450 2.2100 ;
        RECT  5.8250 0.6000 5.9450 0.8400 ;
        RECT  5.0000 1.3200 5.9450 1.4400 ;
        RECT  5.6450 0.7200 5.9450 0.8400 ;
        RECT  5.0000 0.8400 5.7650 0.9600 ;
        RECT  5.0000 1.1750 5.1500 1.4400 ;
        RECT  5.0000 0.7200 5.1200 1.5600 ;
        RECT  4.9850 1.4400 5.1050 2.2100 ;
        RECT  4.9850 0.6000 5.1050 0.8400 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.4050 -0.1800 5.5250 0.6500 ;
        RECT  4.5050 0.4700 4.7450 0.5900 ;
        RECT  4.5050 -0.1800 4.6250 0.5900 ;
        RECT  2.9050 -0.1800 3.0250 0.3800 ;
        RECT  1.4250 -0.1800 1.5450 0.6300 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.4050 1.5600 5.5250 2.7900 ;
        RECT  4.5650 1.7600 4.6850 2.7900 ;
        RECT  3.6650 1.6200 3.9050 2.1500 ;
        RECT  3.6650 1.6200 3.7850 2.7900 ;
        RECT  2.5450 1.9700 2.6650 2.7900 ;
        RECT  1.2650 1.9700 1.3850 2.7900 ;
        RECT  0.1350 1.4600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8250 1.4000 4.6650 1.4000 4.6650 1.6400 4.2650 1.6400 4.2650 2.2100 4.1450 2.2100
                 4.1450 1.5200 4.5450 1.5200 4.5450 0.8300 4.0450 0.8300 4.0450 0.7800 3.8650 0.7800
                 3.8650 0.6600 4.1650 0.6600 4.1650 0.7100 4.6650 0.7100 4.6650 1.1600 4.8250 1.1600 ;
        POLYGON  4.4250 1.4000 3.0850 1.4000 3.0850 2.0900 2.9650 2.0900 2.9650 1.4000 2.4250 1.4000
                 2.4250 1.2800 3.3850 1.2800 3.3850 0.6600 3.5050 0.6600 3.5050 1.2800 4.3050 1.2800
                 4.3050 1.1600 4.4250 1.1600 ;
        POLYGON  4.0450 1.1000 3.8050 1.1000 3.8050 1.0200 3.6250 1.0200 3.6250 0.5400 3.2650 0.5400
                 3.2650 0.6200 2.6650 0.6200 2.6650 0.6000 2.0250 0.6000 2.0250 1.7100 1.7850 1.7100
                 1.7850 1.8200 1.1450 1.8200 1.1450 1.9400 0.9650 1.9400 0.9650 2.0900 0.8450 2.0900
                 0.8450 1.8200 1.0250 1.8200 1.0250 1.7000 1.6650 1.7000 1.6650 1.5900 1.9050 1.5900
                 1.9050 0.8700 1.1100 0.8700 1.1100 0.8400 0.8850 0.8400 0.8850 0.7200 1.2300 0.7200
                 1.2300 0.7500 1.9050 0.7500 1.9050 0.4800 2.3050 0.4800 2.3050 0.3800 2.5450 0.3800
                 2.5450 0.4800 2.7850 0.4800 2.7850 0.5000 3.1450 0.5000 3.1450 0.4200 3.7450 0.4200
                 3.7450 0.9000 3.9250 0.9000 3.9250 0.9800 4.0450 0.9800 ;
        POLYGON  3.1050 1.1600 2.3050 1.1600 2.3050 1.9500 2.0250 1.9500 2.0250 2.0900 1.9050 2.0900
                 1.9050 1.8300 2.1850 1.8300 2.1850 0.8400 2.1450 0.8400 2.1450 0.7200 2.3850 0.7200
                 2.3850 0.8400 2.3050 0.8400 2.3050 1.0400 3.1050 1.0400 ;
        POLYGON  1.7850 1.4500 1.6650 1.4500 1.6650 1.1100 1.0550 1.1100 1.0550 1.1800 0.8150 1.1800
                 0.8150 1.1100 0.6750 1.1100 0.6750 1.5800 0.5550 1.5800 0.5550 0.6800 0.6750 0.6800
                 0.6750 0.9900 1.7850 0.9900 ;
    END
END TLATNCAX3

MACRO TLATNCAX20
    CLASS CORE ;
    FOREIGN TLATNCAX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 15.3700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0600 0.5100 1.5250 ;
        RECT  0.3800 1.0300 0.5000 1.5250 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1350 0.8400 1.5250 ;
        RECT  0.7200 1.1200 0.8400 1.5250 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.6387  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  15.0900 1.2050 15.2100 2.2050 ;
        RECT  15.0100 0.4050 15.1300 1.0300 ;
        RECT  8.1900 1.2050 15.2100 1.3250 ;
        RECT  14.8300 0.9100 15.1300 1.0300 ;
        RECT  14.1700 1.0300 14.9500 1.3250 ;
        RECT  14.2500 1.0300 14.3700 2.2100 ;
        RECT  14.1700 0.4050 14.2900 1.3250 ;
        RECT  13.4100 1.2050 13.5300 2.2100 ;
        RECT  13.1500 0.7900 13.4500 0.9100 ;
        RECT  13.3300 0.4050 13.4500 0.9100 ;
        RECT  12.4900 1.0300 13.2700 1.3250 ;
        RECT  13.1500 0.7900 13.2700 1.3250 ;
        RECT  12.5700 1.0300 12.6900 2.2100 ;
        RECT  12.4900 0.4050 12.6100 1.3250 ;
        RECT  11.7300 1.2050 11.8500 2.2100 ;
        RECT  11.4700 0.7900 11.7700 0.9100 ;
        RECT  11.6500 0.4050 11.7700 0.9100 ;
        RECT  10.8100 1.0300 11.5900 1.3250 ;
        RECT  11.4700 0.7900 11.5900 1.3250 ;
        RECT  10.8900 1.0300 11.0100 2.2100 ;
        RECT  10.8100 0.4050 10.9300 1.3250 ;
        RECT  10.0500 1.2050 10.1700 2.2100 ;
        RECT  9.7900 0.7900 10.0900 0.9100 ;
        RECT  9.9700 0.4050 10.0900 0.9100 ;
        RECT  9.0700 1.0300 9.9100 1.3250 ;
        RECT  9.7900 0.7900 9.9100 1.3250 ;
        RECT  9.2100 1.0300 9.3300 2.2100 ;
        RECT  9.0700 0.4000 9.1900 1.3250 ;
        RECT  8.3700 1.2050 8.4900 2.2100 ;
        RECT  8.2300 1.2050 8.4900 1.4450 ;
        RECT  8.1900 1.1750 8.3500 1.4350 ;
        RECT  8.2300 0.4000 8.3500 1.4450 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 15.3700 0.1800 ;
        RECT  14.5900 -0.1800 14.7100 0.9100 ;
        RECT  13.7500 -0.1800 13.8700 0.9100 ;
        RECT  12.9100 -0.1800 13.0300 0.9100 ;
        RECT  12.0700 -0.1800 12.1900 0.9100 ;
        RECT  11.2300 -0.1800 11.3500 0.9100 ;
        RECT  10.3900 -0.1800 10.5100 0.9100 ;
        RECT  9.5500 -0.1800 9.6700 0.9100 ;
        RECT  8.6500 -0.1800 8.7700 0.9100 ;
        RECT  7.8100 -0.1800 7.9300 0.8700 ;
        RECT  6.2100 0.4600 6.4500 0.5800 ;
        RECT  6.2100 -0.1800 6.3300 0.5800 ;
        RECT  4.7300 0.4600 4.9700 0.5800 ;
        RECT  4.7300 -0.1800 4.8500 0.5800 ;
        RECT  2.9750 -0.1800 3.2150 0.3200 ;
        RECT  2.0150 -0.1800 2.2550 0.3200 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 15.3700 2.7900 ;
        RECT  14.6700 1.4450 14.7900 2.7900 ;
        RECT  13.8300 1.4450 13.9500 2.7900 ;
        RECT  12.9900 1.4450 13.1100 2.7900 ;
        RECT  12.1500 1.4450 12.2700 2.7900 ;
        RECT  11.3100 1.4450 11.4300 2.7900 ;
        RECT  10.4700 1.4450 10.5900 2.7900 ;
        RECT  9.6300 1.4450 9.7500 2.7900 ;
        RECT  8.7900 1.4450 8.9100 2.7900 ;
        RECT  7.9500 1.7100 8.0700 2.7900 ;
        RECT  7.1100 1.7100 7.2300 2.7900 ;
        RECT  6.2700 1.7100 6.3900 2.7900 ;
        RECT  5.4300 1.7100 5.5500 2.7900 ;
        RECT  4.5900 1.7100 4.7100 2.7900 ;
        RECT  3.7500 1.9100 3.8700 2.7900 ;
        RECT  2.9000 2.1500 3.1400 2.2700 ;
        RECT  2.9000 2.1500 3.0200 2.7900 ;
        RECT  1.9400 1.9700 2.1800 2.0900 ;
        RECT  1.9400 1.9700 2.0600 2.7900 ;
        RECT  0.6600 1.6450 0.7800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.0700 1.2300 8.0100 1.2300 8.0100 1.5900 7.6500 1.5900 7.6500 2.2100 7.5300 2.2100
                 7.5300 1.5900 6.8100 1.5900 6.8100 2.2100 6.6900 2.2100 6.6900 1.5900 5.9700 1.5900
                 5.9700 2.2100 5.8500 2.2100 5.8500 1.5900 5.1300 1.5900 5.1300 2.2100 5.0100 2.2100
                 5.0100 1.5900 4.2900 1.5900 4.2900 2.2100 4.1700 2.2100 4.1700 1.4700 7.8900 1.4700
                 7.8900 1.1100 7.1500 1.1100 7.1500 0.8300 7.1100 0.8300 7.1100 0.8200 4.2100 0.8200
                 4.2100 0.7700 4.0900 0.7700 4.0900 0.6500 4.3300 0.6500 4.3300 0.7000 5.3700 0.7000
                 5.3700 0.6500 5.6100 0.6500 5.6100 0.7000 7.1100 0.7000 7.1100 0.5900 7.2300 0.5900
                 7.2300 0.7100 7.2700 0.7100 7.2700 0.9900 8.0700 0.9900 ;
        POLYGON  7.7700 1.3500 4.0500 1.3500 4.0500 1.7900 3.0100 1.7900 3.0100 1.6100 2.4800 1.6100
                 2.4800 1.3700 2.5950 1.3700 2.5950 0.9500 1.7950 0.9500 1.7950 0.8300 2.4950 0.8300
                 2.4950 0.6800 2.7350 0.6800 2.7350 0.8000 2.7150 0.8000 2.7150 1.4900 3.1300 1.4900
                 3.1300 1.6700 3.9300 1.6700 3.9300 1.2300 7.7700 1.2300 ;
        POLYGON  7.0300 1.1100 3.6350 1.1100 3.6350 1.5500 3.3800 1.5500 3.3800 1.4300 3.5150 1.4300
                 3.5150 0.5600 1.6550 0.5600 1.6550 1.0100 1.5350 1.0100 1.5350 0.4400 3.6350 0.4400
                 3.6350 0.9900 7.0300 0.9900 ;
        POLYGON  3.4600 2.0300 2.6450 2.0300 2.6450 1.8500 1.7050 1.8500 1.7050 2.0050 1.5800 2.0050
                 1.5800 2.2250 1.4600 2.2250 1.4600 2.0050 1.0550 2.0050 1.0550 0.9100 0.2400 0.9100
                 0.2400 1.6450 0.3600 1.6450 0.3600 1.8850 0.2400 1.8850 0.2400 1.7650 0.1200 1.7650
                 0.1200 0.6700 0.1350 0.6700 0.1350 0.4300 0.2550 0.4300 0.2550 0.7900 1.0550 0.7900
                 1.0550 0.7500 1.1750 0.7500 1.1750 1.8850 1.5850 1.8850 1.5850 1.7300 2.7650 1.7300
                 2.7650 1.9100 3.4600 1.9100 ;
        POLYGON  2.4750 1.2500 1.4200 1.2500 1.4200 1.7650 1.3000 1.7650 1.3000 1.3700 1.2950 1.3700
                 1.2950 0.4300 1.4150 0.4300 1.4150 1.1300 2.2350 1.1300 2.2350 1.0900 2.4750 1.0900 ;
    END
END TLATNCAX20

MACRO TLATNCAX2
    CLASS CORE ;
    FOREIGN TLATNCAX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.8000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4450 1.0200 0.8000 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        RECT  0.4450 1.0200 0.5650 1.2600 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6550 1.2300 4.9150 1.4500 ;
        RECT  4.6550 1.1800 4.7750 1.5700 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0950 1.1450 1.2150 1.5800 ;
        RECT  0.9400 0.8850 1.1850 1.1450 ;
        RECT  1.0650 0.6800 1.1850 1.2650 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.8000 0.1800 ;
        RECT  4.7350 0.4600 4.9750 0.5800 ;
        RECT  4.7350 -0.1800 4.8550 0.5800 ;
        RECT  3.0550 -0.1800 3.1750 0.3800 ;
        RECT  1.4850 -0.1800 1.6050 0.7300 ;
        RECT  0.6450 -0.1800 0.7650 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.8000 2.7900 ;
        RECT  4.7350 1.6900 4.8550 2.7900 ;
        RECT  3.2550 2.1100 3.3750 2.7900 ;
        RECT  2.2950 2.1200 2.4150 2.7900 ;
        RECT  1.5150 2.1200 1.7550 2.2400 ;
        RECT  1.5150 2.1200 1.6350 2.7900 ;
        RECT  0.6150 1.9400 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.3950 1.7500 5.0950 1.7500 5.0950 1.6300 5.2750 1.6300 5.2750 0.8200 4.4950 0.8200
                 4.4950 0.5200 3.3350 0.5200 3.3350 0.4000 4.6150 0.4000 4.6150 0.7000 5.2750 0.7000
                 5.2750 0.6600 5.3950 0.6600 ;
        POLYGON  5.1550 1.2400 5.0350 1.2400 5.0350 1.0600 4.5350 1.0600 4.5350 1.7100 4.2750 1.7100
                 4.2750 1.7500 4.0350 1.7500 4.0350 1.6300 4.1550 1.6300 4.1550 1.5900 4.4150 1.5900
                 4.4150 1.0600 3.8950 1.0600 3.8950 0.6600 4.0150 0.6600 4.0150 0.9400 5.1550 0.9400 ;
        POLYGON  4.2950 1.4700 4.1750 1.4700 4.1750 1.3500 2.1650 1.3500 2.1650 1.5200 1.9250 1.5200
                 1.9250 1.4000 1.9650 1.4000 1.9650 0.6800 2.0850 0.6800 2.0850 1.2300 3.6350 1.2300
                 3.6350 1.0000 3.7550 1.0000 3.7550 1.2300 4.2950 1.2300 ;
        POLYGON  3.9350 2.2500 3.8150 2.2500 3.8150 1.9900 2.8750 1.9900 2.8750 2.0000 1.0400 2.0000
                 1.0400 1.8200 0.1350 1.8200 0.1350 1.4600 0.1650 1.4600 0.1650 0.6800 0.2850 0.6800
                 0.2850 1.5800 0.2550 1.5800 0.2550 1.7000 1.1600 1.7000 1.1600 1.8800 2.7550 1.8800
                 2.7550 1.8700 3.9350 1.8700 ;
        POLYGON  2.9550 1.7500 2.5700 1.7500 2.5700 1.7600 1.6850 1.7600 1.6850 1.2000 1.3350 1.2000
                 1.3350 1.0800 1.6850 1.0800 1.6850 0.8500 1.7250 0.8500 1.7250 0.4400 2.4750 0.4400
                 2.4750 0.9000 2.3550 0.9000 2.3550 0.5600 1.8450 0.5600 1.8450 0.9700 1.8050 0.9700
                 1.8050 1.6400 2.4500 1.6400 2.4500 1.6300 2.9550 1.6300 ;
    END
END TLATNCAX2

MACRO TLATNCAX16
    CLASS CORE ;
    FOREIGN TLATNCAX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.9200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8450 0.8000 1.1450 ;
        RECT  0.5550 0.9750 0.6750 1.2600 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.8300 1.1750 13.1000 1.4350 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3350 0.7400 6.5750 0.8600 ;
        RECT  5.5550 0.7900 6.4550 0.9100 ;
        RECT  6.0750 1.4900 6.3150 1.6100 ;
        RECT  1.2950 1.3700 6.1950 1.4900 ;
        RECT  5.5550 0.6700 5.6750 1.4900 ;
        RECT  5.2350 1.3700 5.4750 1.6100 ;
        RECT  4.6550 0.7400 4.8950 0.8600 ;
        RECT  4.7100 1.1750 4.8600 1.4900 ;
        RECT  4.3950 1.3700 4.8300 1.6100 ;
        RECT  4.7100 0.7400 4.8300 1.6100 ;
        RECT  3.6950 0.7400 4.0550 0.8600 ;
        RECT  3.4950 1.3700 3.8150 1.6100 ;
        RECT  3.6950 0.7400 3.8150 1.6100 ;
        RECT  2.7950 0.7400 3.2150 0.8600 ;
        RECT  2.6550 1.3700 2.9150 1.6100 ;
        RECT  2.7950 0.7400 2.9150 1.6100 ;
        RECT  1.9550 0.7400 2.3150 0.8600 ;
        RECT  1.8150 1.3700 2.0750 1.6100 ;
        RECT  1.9550 0.7400 2.0750 1.6100 ;
        RECT  0.9750 1.4900 1.4150 1.6100 ;
        RECT  1.2950 0.6800 1.4150 1.6100 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.9200 0.1800 ;
        RECT  13.0700 0.4550 13.3100 0.5750 ;
        RECT  13.1900 -0.1800 13.3100 0.5750 ;
        RECT  11.0950 -0.1800 11.2150 0.4900 ;
        RECT  10.1350 -0.1800 10.2550 0.6700 ;
        RECT  8.4150 0.3700 8.6550 0.4900 ;
        RECT  8.4150 -0.1800 8.5350 0.4900 ;
        RECT  6.8150 -0.1800 6.9350 0.6700 ;
        RECT  5.9750 -0.1800 6.0950 0.6700 ;
        RECT  5.1350 -0.1800 5.2550 0.6700 ;
        RECT  4.2950 -0.1800 4.4150 0.6700 ;
        RECT  3.4550 -0.1800 3.5750 0.6700 ;
        RECT  2.5550 -0.1800 2.6750 0.6650 ;
        RECT  1.7150 -0.1800 1.8350 0.6650 ;
        RECT  0.8750 -0.1800 0.9950 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.9200 2.7900 ;
        RECT  13.0700 1.6350 13.1900 2.7900 ;
        RECT  11.2300 2.0550 11.4700 2.1750 ;
        RECT  11.2300 2.0550 11.3500 2.7900 ;
        RECT  10.3950 2.2300 10.5150 2.7900 ;
        RECT  9.3750 1.9700 9.6150 2.0900 ;
        RECT  9.3750 1.9700 9.4950 2.7900 ;
        RECT  8.4150 1.9700 8.6550 2.0900 ;
        RECT  8.4150 1.9700 8.5350 2.7900 ;
        RECT  7.4550 1.9700 7.6950 2.0900 ;
        RECT  7.4550 1.9700 7.5750 2.7900 ;
        RECT  6.4950 1.9700 6.7350 2.1100 ;
        RECT  6.4950 1.9700 6.6150 2.7900 ;
        RECT  5.6550 1.9700 5.8950 2.1100 ;
        RECT  5.6550 1.9700 5.7750 2.7900 ;
        RECT  4.8150 1.9700 5.0550 2.1100 ;
        RECT  4.8150 1.9700 4.9350 2.7900 ;
        RECT  3.9150 1.9700 4.1550 2.1150 ;
        RECT  3.9150 1.9700 4.0350 2.7900 ;
        RECT  3.0750 1.9700 3.3150 2.1150 ;
        RECT  3.0750 1.9700 3.1950 2.7900 ;
        RECT  2.2350 1.9700 2.4750 2.1150 ;
        RECT  2.2350 1.9700 2.3550 2.7900 ;
        RECT  1.3950 1.9700 1.6350 2.1150 ;
        RECT  1.3950 1.9700 1.5150 2.7900 ;
        RECT  0.5550 1.9700 0.7950 2.1150 ;
        RECT  0.5550 1.9700 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.7300 1.6350 13.6100 1.6350 13.6100 1.7550 13.4900 1.7550 13.4900 1.5150
                 13.6100 1.5150 13.6100 0.8150 12.8300 0.8150 12.8300 0.5000 11.7700 0.5000
                 11.7700 0.7300 10.8550 0.7300 10.8550 0.5000 10.4950 0.5000 10.4950 0.9700
                 9.2750 0.9700 9.2750 1.1200 9.0350 1.1200 9.0350 0.9700 8.0350 0.9700 8.0350 1.1200
                 7.7950 1.1200 7.7950 0.8500 10.3750 0.8500 10.3750 0.3800 10.9750 0.3800
                 10.9750 0.6100 11.6500 0.6100 11.6500 0.3800 12.0100 0.3800 12.0100 0.3600
                 12.2500 0.3600 12.2500 0.3800 12.9500 0.3800 12.9500 0.6950 13.6100 0.6950
                 13.6100 0.6200 13.7300 0.6200 ;
        POLYGON  13.3500 1.2000 13.2300 1.2000 13.2300 1.0550 12.7100 1.0550 12.7100 1.9350
                 9.9400 1.9350 9.9400 1.8500 0.1350 1.8500 0.1350 1.4300 0.3150 1.4300 0.3150 0.6800
                 0.4350 0.6800 0.4350 1.5500 0.2550 1.5500 0.2550 1.7300 10.0600 1.7300 10.0600 1.8150
                 12.5900 1.8150 12.5900 1.4150 11.8700 1.4150 11.8700 1.1750 11.9900 1.1750
                 11.9900 1.2950 12.5900 1.2950 12.5900 0.9350 13.3500 0.9350 ;
        POLYGON  12.4700 0.9700 11.7500 0.9700 11.7500 1.5350 12.0500 1.5350 12.0500 1.5750
                 12.1700 1.5750 12.1700 1.6950 11.9300 1.6950 11.9300 1.6550 11.6300 1.6550
                 11.6300 1.4200 11.0500 1.4200 11.0500 1.0900 11.1700 1.0900 11.1700 1.3000
                 11.6300 1.3000 11.6300 0.8500 12.3500 0.8500 12.3500 0.6200 12.4700 0.6200 ;
        POLYGON  11.5100 1.1800 11.3900 1.1800 11.3900 0.9700 10.7350 0.9700 10.7350 1.3600
                 10.9300 1.3600 10.9300 1.6950 10.8100 1.6950 10.8100 1.4800 10.6150 1.4800
                 10.6150 1.3600 6.9550 1.3600 6.9550 1.1100 7.0750 1.1100 7.0750 1.2400 8.2550 1.2400
                 8.2550 1.0900 8.3750 1.0900 8.3750 1.2400 10.1150 1.2400 10.1150 1.1100 10.2350 1.1100
                 10.2350 1.2400 10.6150 1.2400 10.6150 0.6200 10.7350 0.6200 10.7350 0.8500
                 11.5100 0.8500 ;
        POLYGON  10.0950 1.6100 9.8550 1.6100 9.8550 1.6000 9.1350 1.6000 9.1350 1.6100 8.8950 1.6100
                 8.8950 1.6000 8.1750 1.6000 8.1750 1.6100 7.9350 1.6100 7.9350 1.6000 7.2150 1.6000
                 7.2150 1.6100 6.9750 1.6100 6.9750 1.6000 6.7150 1.6000 6.7150 1.1800 6.1950 1.1800
                 6.1950 1.0600 6.7150 1.0600 6.7150 0.8600 7.4600 0.8600 7.4600 0.6100 9.5550 0.6100
                 9.5550 0.7300 7.5800 0.7300 7.5800 0.9800 6.8350 0.9800 6.8350 1.4800 9.9750 1.4800
                 9.9750 1.4900 10.0950 1.4900 ;
    END
END TLATNCAX16

MACRO TLATNCAX12
    CLASS CORE ;
    FOREIGN TLATNCAX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.7300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2300 0.8550 1.3800 ;
        RECT  0.5950 1.0800 0.7150 1.3800 ;
        RECT  0.3550 1.0800 0.7150 1.2000 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.9300 1.4650 10.0800 1.7250 ;
        RECT  9.9300 1.3400 10.0500 1.7250 ;
        RECT  9.8950 1.2200 10.0150 1.4600 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2750 1.4000 4.5150 1.5800 ;
        RECT  1.2150 0.8400 4.5150 0.9600 ;
        RECT  4.3950 0.4000 4.5150 0.9600 ;
        RECT  1.2150 1.3200 4.3950 1.4400 ;
        RECT  3.4350 1.3200 3.6750 1.5800 ;
        RECT  3.5550 0.4000 3.6750 0.9600 ;
        RECT  2.5950 1.3200 2.8350 1.5800 ;
        RECT  2.7150 0.4000 2.8350 0.9600 ;
        RECT  1.7550 1.3200 1.9950 1.5800 ;
        RECT  1.8750 0.4000 1.9950 0.9600 ;
        RECT  1.2150 1.1750 1.3800 1.4400 ;
        RECT  0.9750 1.3400 1.3350 1.4600 ;
        RECT  1.2150 0.8000 1.3350 1.4600 ;
        RECT  1.0350 0.8000 1.3350 0.9200 ;
        RECT  1.0350 0.4000 1.1550 0.9200 ;
        RECT  0.9750 1.3400 1.0950 1.5800 ;
        END
    END ECK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.7300 0.1800 ;
        RECT  9.9750 0.5000 10.2150 0.6200 ;
        RECT  10.0950 -0.1800 10.2150 0.6200 ;
        RECT  8.0750 -0.1800 8.1950 0.7300 ;
        RECT  6.4150 0.5500 6.6550 0.6700 ;
        RECT  6.4150 -0.1800 6.5350 0.6700 ;
        RECT  4.8150 -0.1800 4.9350 0.9150 ;
        RECT  3.9750 -0.1800 4.0950 0.7200 ;
        RECT  3.1350 -0.1800 3.2550 0.7200 ;
        RECT  2.2950 -0.1800 2.4150 0.7200 ;
        RECT  1.4550 -0.1800 1.5750 0.7200 ;
        RECT  0.6150 -0.1800 0.7350 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.7300 2.7900 ;
        RECT  10.0550 1.8450 10.1750 2.7900 ;
        RECT  8.3350 2.2000 8.4550 2.7900 ;
        RECT  7.3150 2.1000 7.5550 2.2200 ;
        RECT  7.3150 2.1000 7.4350 2.7900 ;
        RECT  6.3550 2.1000 6.5950 2.2200 ;
        RECT  6.3550 2.1000 6.4750 2.7900 ;
        RECT  5.3950 2.1200 5.6350 2.2400 ;
        RECT  5.3950 2.1200 5.5150 2.7900 ;
        RECT  4.7550 2.1200 4.9950 2.2400 ;
        RECT  4.7550 2.1200 4.8750 2.7900 ;
        RECT  3.8550 1.9400 4.0950 2.0600 ;
        RECT  3.8550 1.9400 3.9750 2.7900 ;
        RECT  3.0150 1.9400 3.2550 2.0600 ;
        RECT  3.0150 1.9400 3.1350 2.7900 ;
        RECT  2.1750 1.9400 2.4150 2.0600 ;
        RECT  2.1750 1.9400 2.2950 2.7900 ;
        RECT  1.3350 1.9400 1.5750 2.0600 ;
        RECT  1.3350 1.9400 1.4550 2.7900 ;
        RECT  0.4950 1.9800 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.5950 2.2100 10.4750 2.2100 10.4750 1.6800 10.4550 1.6800 10.4550 0.8600
                 9.7350 0.8600 9.7350 0.5700 8.4350 0.5700 8.4350 1.1600 8.3150 1.1600 8.3150 1.1800
                 8.0750 1.1800 8.0750 1.1600 6.9150 1.1600 6.9150 1.2000 6.6750 1.2000 6.6750 1.0400
                 8.3150 1.0400 8.3150 0.4500 9.8550 0.4500 9.8550 0.7400 10.4550 0.7400 10.4550 0.6300
                 10.5750 0.6300 10.5750 1.5600 10.5950 1.5600 ;
        POLYGON  10.3350 1.2200 10.2150 1.2200 10.2150 1.1000 9.7750 1.1000 9.7750 1.7000 9.5350 1.7000
                 9.5350 1.7400 9.2950 1.7400 9.2950 1.6200 9.4150 1.6200 9.4150 1.5800 9.6550 1.5800
                 9.6550 1.1000 9.1150 1.1000 9.1150 0.8100 8.9750 0.8100 8.9750 0.6900 9.2350 0.6900
                 9.2350 0.9800 10.3350 0.9800 ;
        POLYGON  9.5350 1.4600 9.4150 1.4600 9.4150 1.4400 5.4150 1.4400 5.4150 1.5200 5.1150 1.5200
                 5.1150 1.4000 5.2950 1.4000 5.2950 0.6750 5.4150 0.6750 5.4150 1.3200 5.5950 1.3200
                 5.5950 1.3000 5.8350 1.3000 5.8350 1.3200 7.0350 1.3200 7.0350 1.2800 7.2750 1.2800
                 7.2750 1.3200 8.8750 1.3200 8.8750 0.9700 8.9950 0.9700 8.9950 1.3200 9.4150 1.3200
                 9.4150 1.2200 9.5350 1.2200 ;
        POLYGON  9.1950 2.2400 9.0750 2.2400 9.0750 2.1200 9.0300 2.1200 9.0300 2.0800 8.2350 2.0800
                 8.2350 1.9800 6.2350 1.9800 6.2350 2.0000 4.5450 2.0000 4.5450 1.8200 0.1350 1.8200
                 0.1350 1.5800 0.1150 1.5800 0.1150 0.8000 0.1350 0.8000 0.1350 0.6800 0.2550 0.6800
                 0.2550 0.9200 0.2350 0.9200 0.2350 1.4600 0.2550 1.4600 0.2550 1.7000 4.6650 1.7000
                 4.6650 1.8800 6.1150 1.8800 6.1150 1.8600 8.3550 1.8600 8.3550 1.9600 9.1500 1.9600
                 9.1500 2.0000 9.1950 2.0000 ;
        POLYGON  8.0350 1.7400 5.7500 1.7400 5.7500 1.7600 4.8750 1.7600 4.8750 1.2000 4.1950 1.2000
                 4.1950 1.0800 5.0550 1.0800 5.0550 0.4350 5.7050 0.4350 5.7050 0.5500 5.9500 0.5500
                 5.9500 0.7900 6.8900 0.7900 6.8900 0.7400 7.3950 0.7400 7.3950 0.8600 7.0100 0.8600
                 7.0100 0.9100 5.8300 0.9100 5.8300 0.6700 5.5850 0.6700 5.5850 0.5550 5.1750 0.5550
                 5.1750 1.2000 4.9950 1.2000 4.9950 1.6400 5.6300 1.6400 5.6300 1.6200 8.0350 1.6200 ;
    END
END TLATNCAX12

MACRO TIELO
    CLASS CORE ;
    FOREIGN TIELO 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.8700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1204  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.5450 0.2550 0.9600 ;
        RECT  0.1350 0.5300 0.2550 0.9600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.8700 0.1800 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.8700 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  0.4550 1.2000 0.2550 1.2000 0.2550 1.9900 0.1350 1.9900 0.1350 1.0800 0.4550 1.0800 ;
    END
END TIELO

MACRO TIEHI
    CLASS CORE ;
    FOREIGN TIEHI 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.8700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1820  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 1.3800 0.2550 2.0300 ;
        RECT  0.0700 1.4650 0.2550 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.8700 0.1800 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.8700 2.7900 ;
        RECT  0.5550 1.3800 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  0.4150 1.2600 0.2950 1.2600 0.2950 0.9200 0.1350 0.9200 0.1350 0.6800 0.2550 0.6800
                 0.2550 0.8000 0.4150 0.8000 ;
    END
END TIEHI

MACRO TBUFXL
    CLASS CORE ;
    FOREIGN TBUFXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4350 1.1600 1.4150 1.2800 ;
        RECT  0.4350 1.0250 0.8000 1.2800 ;
        RECT  0.6500 0.8850 0.8000 1.2800 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2200 0.3600 2.7250 0.4800 ;
        RECT  1.2150 0.4400 2.3400 0.5600 ;
        RECT  0.8150 1.4000 1.6550 1.5200 ;
        RECT  1.5350 0.9200 1.6550 1.5200 ;
        RECT  1.2150 0.9200 1.6550 1.0400 ;
        RECT  1.1750 1.4000 1.4350 1.6700 ;
        RECT  1.2150 0.4400 1.3350 1.0400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2450 0.7600 3.3650 1.6050 ;
        RECT  2.9700 1.4650 3.3450 1.7250 ;
        RECT  3.2250 0.6400 3.3450 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.8450 -0.1800 2.9650 0.7600 ;
        RECT  2.8050 0.6400 2.9250 0.8800 ;
        RECT  1.8450 -0.1800 2.0850 0.3200 ;
        RECT  0.9750 -0.1800 1.0950 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.7450 2.0850 2.8650 2.7900 ;
        RECT  1.0350 2.2900 1.2750 2.7900 ;
        RECT  0.1350 1.8800 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1850 2.1850 3.0650 2.1850 3.0650 1.9650 2.3900 1.9650 2.3900 2.1700 1.2100 2.1700
                 1.2100 2.1100 0.6150 2.1100 0.6150 1.7600 0.1950 1.7600 0.1950 0.7850 0.2750 0.7850
                 0.2750 0.6200 0.3950 0.6200 0.3950 0.9050 0.3150 0.9050 0.3150 1.6400 0.7350 1.6400
                 0.7350 1.9900 1.3300 1.9900 1.3300 2.0500 2.2700 2.0500 2.2700 1.8450 3.1850 1.8450 ;
        POLYGON  3.1250 1.1400 2.5250 1.1400 2.5250 1.4850 2.1650 1.4850 2.1650 1.7250 2.0450 1.7250
                 2.0450 1.3650 2.4050 1.3650 2.4050 0.8200 2.3250 0.8200 2.3250 0.7000 2.5650 0.7000
                 2.5650 0.8200 2.5250 0.8200 2.5250 1.0200 3.1250 1.0200 ;
        POLYGON  2.2850 1.2450 1.8950 1.2450 1.8950 1.9300 1.5150 1.9300 1.5150 1.8100 1.7750 1.8100
                 1.7750 0.8000 1.4550 0.8000 1.4550 0.6800 1.8950 0.6800 1.8950 1.1250 2.2850 1.1250 ;
    END
END TBUFXL

MACRO TBUFX8
    CLASS CORE ;
    FOREIGN TBUFX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2760  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3150 0.9400 2.4350 1.1800 ;
        RECT  0.6500 0.9900 2.4350 1.1100 ;
        RECT  1.5550 0.9900 1.7950 1.1400 ;
        RECT  0.3350 1.3150 0.8000 1.4350 ;
        RECT  0.6500 0.9900 0.8000 1.4350 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6150 0.3600 5.8550 0.4800 ;
        RECT  3.4350 0.4900 5.7350 0.6100 ;
        RECT  5.6150 0.3600 5.7350 0.6100 ;
        RECT  4.3950 0.3650 4.6350 0.6100 ;
        RECT  3.6750 0.3650 3.9150 0.6100 ;
        RECT  2.5550 0.4400 3.5550 0.5600 ;
        RECT  1.0950 1.3400 2.6750 1.4600 ;
        RECT  2.5550 0.4400 2.6750 1.4600 ;
        RECT  1.1750 1.2300 1.4350 1.4600 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2150 0.8400 9.0150 0.9600 ;
        RECT  8.8950 0.6700 9.0150 0.9600 ;
        RECT  8.7550 0.8400 8.8750 2.2100 ;
        RECT  6.7400 1.3200 8.8750 1.4400 ;
        RECT  8.0550 0.6700 8.1750 0.9600 ;
        RECT  7.9150 1.3200 8.0350 2.2100 ;
        RECT  7.2150 0.6700 7.3350 0.9600 ;
        RECT  7.0750 1.3200 7.1950 2.2100 ;
        RECT  6.7400 1.1750 6.8900 1.4400 ;
        RECT  6.2350 1.5900 6.8600 1.7100 ;
        RECT  6.7400 0.9900 6.8600 1.7100 ;
        RECT  6.3750 0.9900 6.8600 1.1100 ;
        RECT  6.3750 0.6700 6.4950 1.1100 ;
        RECT  6.2350 1.5900 6.3550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  9.3150 -0.1800 9.4350 0.7200 ;
        RECT  8.4750 -0.1800 8.5950 0.7200 ;
        RECT  7.6350 -0.1800 7.7550 0.7200 ;
        RECT  6.7950 -0.1800 6.9150 0.7200 ;
        RECT  5.8950 0.6800 6.1350 0.8000 ;
        RECT  5.9750 -0.1800 6.0950 0.8000 ;
        RECT  4.9950 -0.1800 5.2350 0.3700 ;
        RECT  4.0350 -0.1800 4.2750 0.3700 ;
        RECT  3.0750 -0.1800 3.3150 0.3200 ;
        RECT  2.2350 -0.1800 2.3550 0.8100 ;
        RECT  0.7750 0.5100 1.0150 0.6300 ;
        RECT  0.7750 -0.1800 0.8950 0.6300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  9.1750 1.5600 9.2950 2.7900 ;
        RECT  8.3350 1.5600 8.4550 2.7900 ;
        RECT  7.4950 1.5600 7.6150 2.7900 ;
        RECT  6.6550 1.8300 6.7750 2.7900 ;
        RECT  5.8150 1.5900 5.9350 2.7900 ;
        RECT  4.4150 2.0250 4.6550 2.1450 ;
        RECT  4.4150 2.0250 4.5350 2.7900 ;
        RECT  2.7150 2.2400 2.9550 2.7900 ;
        RECT  1.8750 1.8950 1.9950 2.7900 ;
        RECT  1.0350 1.8950 1.1550 2.7900 ;
        RECT  0.1350 1.8900 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.5750 1.4700 5.6950 1.4700 5.6950 2.1950 4.7750 2.1950 4.7750 1.9050 4.2700 1.9050
                 4.2700 2.1950 3.0900 2.1950 3.0900 2.1200 2.2950 2.1200 2.2950 1.7600 1.5750 1.7600
                 1.5750 1.9400 1.4550 1.9400 1.4550 1.7600 0.6750 1.7600 0.6750 1.9400 0.5550 1.9400
                 0.5550 1.7600 0.0950 1.7600 0.0950 0.7350 0.1350 0.7350 0.1350 0.6150 0.2550 0.6150
                 0.2550 0.7350 0.5200 0.7350 0.5200 0.7500 1.1950 0.7500 1.1950 0.6800 1.7750 0.6800
                 1.7750 0.8000 1.3150 0.8000 1.3150 0.8700 0.4000 0.8700 0.4000 0.8550 0.2150 0.8550
                 0.2150 1.6400 2.4150 1.6400 2.4150 2.0000 3.2100 2.0000 3.2100 2.0750 4.1500 2.0750
                 4.1500 1.7850 4.8950 1.7850 4.8950 2.0750 5.5750 2.0750 5.5750 1.3500 6.4550 1.3500
                 6.4550 1.2300 6.5750 1.2300 ;
        POLYGON  6.2150 1.2300 6.0950 1.2300 6.0950 1.0400 5.3750 1.0400 5.3750 1.9550 5.0550 1.9550
                 5.0550 1.8350 5.2550 1.8350 5.2550 1.6650 4.0150 1.6650 4.0150 1.9550 3.7750 1.9550
                 3.7750 1.8350 3.8950 1.8350 3.8950 1.5450 5.2550 1.5450 5.2550 1.0400 3.6750 1.0400
                 3.6750 0.8500 3.5550 0.8500 3.5550 0.7300 3.7950 0.7300 3.7950 0.9200 4.5150 0.9200
                 4.5150 0.7300 4.7550 0.7300 4.7550 0.9200 5.4750 0.9200 5.4750 0.7300 5.7150 0.7300
                 5.7150 0.9200 6.2150 0.9200 ;
        POLYGON  5.1350 1.2800 3.3150 1.2800 3.3150 1.7600 3.4350 1.7600 3.4350 1.8800 3.1950 1.8800
                 3.1950 0.8000 2.7950 0.8000 2.7950 0.6800 3.3150 0.6800 3.3150 1.1600 5.1350 1.1600 ;
    END
END TBUFX8

MACRO TBUFX6
    CLASS CORE ;
    FOREIGN TBUFX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2760  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3150 0.9400 2.4350 1.1800 ;
        RECT  0.6500 0.9900 2.4350 1.1100 ;
        RECT  1.5550 0.9900 1.7950 1.1400 ;
        RECT  0.3350 1.3150 0.8000 1.4350 ;
        RECT  0.6500 0.9900 0.8000 1.4350 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7200 0.3600 5.9600 0.4800 ;
        RECT  3.5150 0.4900 5.8400 0.6100 ;
        RECT  5.7200 0.3600 5.8400 0.6100 ;
        RECT  4.5000 0.3650 4.7400 0.6100 ;
        RECT  3.7800 0.3650 4.0200 0.6100 ;
        RECT  2.5550 0.4400 3.6350 0.5600 ;
        RECT  1.0950 1.3400 2.6750 1.4600 ;
        RECT  2.5550 0.4400 2.6750 1.4600 ;
        RECT  1.1750 1.2300 1.4350 1.4600 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0368  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3200 0.8400 8.2800 0.9600 ;
        RECT  8.1600 0.6700 8.2800 0.9600 ;
        RECT  8.1400 0.8400 8.2600 2.2100 ;
        RECT  6.7400 1.3200 8.2600 1.4400 ;
        RECT  7.3200 0.6700 7.4400 0.9600 ;
        RECT  7.3000 1.3200 7.4200 2.2100 ;
        RECT  6.7400 1.1750 6.8900 1.4400 ;
        RECT  6.4600 1.5900 6.8600 1.7100 ;
        RECT  6.7400 0.9900 6.8600 1.7100 ;
        RECT  6.4800 0.9900 6.8600 1.1100 ;
        RECT  6.4800 0.6700 6.6000 1.1100 ;
        RECT  6.4600 1.5900 6.5800 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.5800 -0.1800 8.7000 0.7200 ;
        RECT  7.7400 -0.1800 7.8600 0.7200 ;
        RECT  6.9000 -0.1800 7.0200 0.7200 ;
        RECT  6.0000 0.6800 6.2400 0.8000 ;
        RECT  6.0800 -0.1800 6.2000 0.8000 ;
        RECT  5.1000 -0.1800 5.3400 0.3700 ;
        RECT  4.1400 -0.1800 4.3800 0.3700 ;
        RECT  3.1800 -0.1800 3.4200 0.3200 ;
        RECT  2.2350 -0.1800 2.3550 0.8100 ;
        RECT  0.7750 0.5100 1.0150 0.6300 ;
        RECT  0.7750 -0.1800 0.8950 0.6300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.5600 1.5600 8.6800 2.7900 ;
        RECT  7.7200 1.5600 7.8400 2.7900 ;
        RECT  6.8800 1.8300 7.0000 2.7900 ;
        RECT  6.0400 1.5900 6.1600 2.7900 ;
        RECT  4.6400 2.0250 4.8800 2.1450 ;
        RECT  4.6400 2.0250 4.7600 2.7900 ;
        RECT  2.7150 2.2400 2.9550 2.7900 ;
        RECT  1.8750 1.8950 1.9950 2.7900 ;
        RECT  1.0350 1.8950 1.1550 2.7900 ;
        RECT  0.1350 1.8900 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.6200 1.4700 5.8250 1.4700 5.8250 2.1950 5.0000 2.1950 5.0000 1.9050 4.5200 1.9050
                 4.5200 2.1950 3.6200 2.1950 3.6200 2.1200 2.2950 2.1200 2.2950 1.7600 1.5750 1.7600
                 1.5750 1.9400 1.4550 1.9400 1.4550 1.7600 0.6750 1.7600 0.6750 1.9400 0.5550 1.9400
                 0.5550 1.7600 0.0950 1.7600 0.0950 0.7350 0.1350 0.7350 0.1350 0.6150 0.2550 0.6150
                 0.2550 0.7350 0.5200 0.7350 0.5200 0.7500 1.1950 0.7500 1.1950 0.6800 1.7750 0.6800
                 1.7750 0.8000 1.3150 0.8000 1.3150 0.8700 0.4000 0.8700 0.4000 0.8550 0.2150 0.8550
                 0.2150 1.6400 2.4150 1.6400 2.4150 2.0000 3.7400 2.0000 3.7400 2.0750 4.4000 2.0750
                 4.4000 1.7850 5.1200 1.7850 5.1200 2.0750 5.7050 2.0750 5.7050 1.3500 6.5000 1.3500
                 6.5000 1.2300 6.6200 1.2300 ;
        POLYGON  6.2600 1.2300 6.1400 1.2300 6.1400 1.0400 5.5000 1.0400 5.5000 1.8350 5.5200 1.8350
                 5.5200 1.9550 5.2800 1.9550 5.2800 1.8350 5.3800 1.8350 5.3800 1.6650 4.2800 1.6650
                 4.2800 1.9550 3.9600 1.9550 3.9600 1.8350 4.1600 1.8350 4.1600 1.5450 5.3800 1.5450
                 5.3800 1.0400 3.7800 1.0400 3.7800 0.8500 3.6600 0.8500 3.6600 0.7300 3.9000 0.7300
                 3.9000 0.9200 4.6200 0.9200 4.6200 0.7300 4.8600 0.7300 4.8600 0.9200 5.5800 0.9200
                 5.5800 0.7300 5.8200 0.7300 5.8200 0.9200 6.2600 0.9200 ;
        POLYGON  5.2600 1.2800 3.3950 1.2800 3.3950 1.7600 3.4350 1.7600 3.4350 1.8800 3.1950 1.8800
                 3.1950 1.7600 3.2750 1.7600 3.2750 0.8000 2.7950 0.8000 2.7950 0.6800 3.3950 0.6800
                 3.3950 1.1600 5.2600 1.1600 ;
    END
END TBUFX6

MACRO TBUFX4
    CLASS CORE ;
    FOREIGN TBUFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3000 1.0400 1.1400 1.1600 ;
        RECT  0.3600 0.8850 0.5100 1.1600 ;
        RECT  0.3000 1.0000 0.4200 1.2400 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5550 0.9900 2.8350 1.1100 ;
        RECT  2.7150 0.4100 2.8350 1.1100 ;
        RECT  2.0750 0.4100 2.8350 0.5300 ;
        RECT  1.2600 0.4800 2.1950 0.6000 ;
        RECT  1.2600 1.2300 1.7250 1.3800 ;
        RECT  0.5600 1.2800 1.5850 1.4000 ;
        RECT  1.2600 0.4800 1.3800 1.4000 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2550 1.3150 4.3750 2.2100 ;
        RECT  3.5350 0.7600 4.3350 0.8800 ;
        RECT  4.2150 0.5900 4.3350 0.8800 ;
        RECT  3.5350 1.3150 4.3750 1.4350 ;
        RECT  3.5350 1.1750 3.7000 1.4350 ;
        RECT  3.5350 0.7100 3.6550 1.8300 ;
        RECT  3.4150 1.7100 3.5350 2.2100 ;
        RECT  3.3750 0.7100 3.6550 0.8300 ;
        RECT  3.3750 0.5900 3.4950 0.8300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  4.6350 -0.1800 4.7550 0.6400 ;
        RECT  3.7950 -0.1800 3.9150 0.6400 ;
        RECT  2.9550 -0.1800 3.0750 0.6400 ;
        RECT  1.7150 -0.1800 1.9550 0.3600 ;
        RECT  0.7800 -0.1800 0.9000 0.7100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  4.6750 1.5600 4.7950 2.7900 ;
        RECT  3.7750 1.6200 4.0150 2.1500 ;
        RECT  3.7750 1.6200 3.8950 2.7900 ;
        RECT  2.9150 1.7100 3.0350 2.7900 ;
        RECT  0.9750 2.1000 1.2150 2.2200 ;
        RECT  0.9750 2.1000 1.0950 2.7900 ;
        RECT  0.1350 1.7600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.4150 1.5900 2.7950 1.5900 2.7950 1.8000 2.5300 1.8000 2.5300 2.2500 1.6150 2.2500
                 1.6150 1.9800 0.6750 1.9800 0.6750 2.2100 0.5550 2.2100 0.5550 1.6400 0.0600 1.6400
                 0.0600 0.6450 0.1400 0.6450 0.1400 0.5250 0.2600 0.5250 0.2600 0.7650 0.1800 0.7650
                 0.1800 1.5200 0.6750 1.5200 0.6750 1.8600 1.7350 1.8600 1.7350 2.1300 2.4100 2.1300
                 2.4100 1.6800 2.6750 1.6800 2.6750 1.4700 3.2950 1.4700 3.2950 1.2200 3.4150 1.2200 ;
        POLYGON  3.0750 1.3500 2.4350 1.3500 2.4350 1.5600 2.2550 1.5600 2.2550 2.0100 2.1350 2.0100
                 2.1350 1.4400 2.3150 1.4400 2.3150 0.6500 2.5950 0.6500 2.5950 0.7700 2.4350 0.7700
                 2.4350 1.2300 2.9550 1.2300 2.9550 0.9100 3.0750 0.9100 ;
        POLYGON  2.1950 1.3200 1.9650 1.3200 1.9650 1.7400 1.4550 1.7400 1.4550 1.6200 1.8450 1.6200
                 1.8450 0.8400 1.5000 0.8400 1.5000 0.7200 1.9650 0.7200 1.9650 1.2000 2.1950 1.2000 ;
    END
END TBUFX4

MACRO TBUFX3
    CLASS CORE ;
    FOREIGN TBUFX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0000 1.2900 1.1200 ;
        RECT  0.3900 0.8850 0.5100 1.2400 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.8450 0.9600 3.0000 1.2000 ;
        RECT  2.8800 0.4400 3.0000 1.2000 ;
        RECT  1.4100 0.4400 3.0000 0.5600 ;
        RECT  1.4650 1.2300 1.7250 1.3800 ;
        RECT  1.4100 0.4400 1.5300 1.3600 ;
        RECT  0.7100 1.2400 1.7250 1.3600 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3850 1.5600 4.5050 2.2100 ;
        RECT  4.3800 0.6200 4.5000 0.8600 ;
        RECT  3.8400 1.5600 4.5050 1.6800 ;
        RECT  4.2000 0.7400 4.5000 0.8600 ;
        RECT  3.8400 0.8600 4.3200 0.9800 ;
        RECT  3.8400 1.4650 3.9900 1.7250 ;
        RECT  3.4250 1.8000 3.9600 1.9200 ;
        RECT  3.8400 0.7900 3.9600 1.9200 ;
        RECT  3.5400 0.7900 3.9600 0.9100 ;
        RECT  3.5400 0.6200 3.6600 0.9100 ;
        RECT  3.4250 1.8000 3.5450 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  3.9600 -0.1800 4.0800 0.6700 ;
        RECT  3.1200 -0.1800 3.2400 0.6700 ;
        RECT  2.0400 -0.1800 2.2800 0.3200 ;
        RECT  0.9300 -0.1800 1.0500 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  3.9050 2.0400 4.0250 2.7900 ;
        RECT  3.0050 1.8000 3.1250 2.7900 ;
        RECT  0.9750 2.1000 1.2150 2.2200 ;
        RECT  0.9750 2.1000 1.0950 2.7900 ;
        RECT  0.1350 1.7200 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.7200 1.6800 2.8850 1.6800 2.8850 1.8000 2.7250 1.8000 2.7250 2.2500 2.0750 2.2500
                 2.0750 1.9800 0.6750 1.9800 0.6750 2.2100 0.5550 2.2100 0.5550 1.6000 0.1200 1.6000
                 0.1200 0.6450 0.2900 0.6450 0.2900 0.5250 0.4100 0.5250 0.4100 0.7650 0.2400 0.7650
                 0.2400 1.4800 0.6750 1.4800 0.6750 1.8600 2.1950 1.8600 2.1950 2.1300 2.6050 2.1300
                 2.6050 1.6800 2.7650 1.6800 2.7650 1.5600 3.6000 1.5600 3.6000 1.2200 3.7200 1.2200 ;
        POLYGON  3.3800 1.4400 2.6450 1.4400 2.6450 1.5600 2.4850 1.5600 2.4850 2.0100 2.3650 2.0100
                 2.3650 1.4400 2.5250 1.4400 2.5250 0.8000 2.5200 0.8000 2.5200 0.6800 2.7600 0.6800
                 2.7600 0.8000 2.6450 0.8000 2.6450 1.3200 3.2600 1.3200 3.2600 0.9400 3.3800 0.9400 ;
        POLYGON  2.4050 1.3200 1.9650 1.3200 1.9650 1.6200 1.6950 1.6200 1.6950 1.7400 1.4550 1.7400
                 1.4550 1.6200 1.5750 1.6200 1.5750 1.5000 1.8450 1.5000 1.8450 0.8000 1.6500 0.8000
                 1.6500 0.6800 1.9650 0.6800 1.9650 1.2000 2.4050 1.2000 ;
    END
END TBUFX3

MACRO TBUFX20
    CLASS CORE ;
    FOREIGN TBUFX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 19.7200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.0800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0850 0.9400 10.8650 1.0600 ;
        RECT  6.0850 0.7600 6.2050 1.0600 ;
        RECT  5.6650 0.7600 6.2050 0.8800 ;
        RECT  5.6650 0.4100 5.7850 0.8800 ;
        RECT  5.0650 0.4100 5.7850 0.5300 ;
        RECT  4.5850 0.7850 5.1850 0.9050 ;
        RECT  5.0650 0.4100 5.1850 0.9050 ;
        RECT  4.8650 0.7850 4.9850 1.1500 ;
        RECT  4.5850 0.3600 4.7050 0.9050 ;
        RECT  3.8850 0.3600 4.7050 0.4800 ;
        RECT  2.9450 0.7800 4.0050 0.9000 ;
        RECT  3.8850 0.3600 4.0050 0.9000 ;
        RECT  3.3850 0.7800 3.5050 1.1000 ;
        RECT  2.9450 0.3600 3.0650 0.9000 ;
        RECT  2.0850 0.3600 3.0650 0.4800 ;
        RECT  1.6050 0.7800 2.2050 0.9000 ;
        RECT  2.0850 0.3600 2.2050 0.9000 ;
        RECT  2.0250 0.7800 2.1450 1.1200 ;
        RECT  1.6250 0.7800 1.7450 1.1200 ;
        RECT  1.6050 0.3600 1.7250 0.9000 ;
        RECT  0.6050 0.3600 1.7250 0.4800 ;
        RECT  0.3050 0.9400 0.7250 1.0600 ;
        RECT  0.6050 0.3600 0.7250 1.0600 ;
        RECT  0.3050 0.9400 0.5650 1.0900 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3926  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.7560  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.5193  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.8450 1.2200 4.2250 1.3400 ;
        RECT  4.1050 1.0700 4.2250 1.3400 ;
        RECT  2.9150 1.2200 3.1750 1.3800 ;
        RECT  2.8450 1.0700 2.9650 1.3400 ;
        END
    END OE
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.4560  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  19.0450 1.4000 19.1650 2.1700 ;
        RECT  17.2450 0.7600 19.0450 0.8800 ;
        RECT  18.9250 0.5900 19.0450 0.8800 ;
        RECT  18.8650 1.4000 19.1650 1.5200 ;
        RECT  11.6650 1.2800 18.9850 1.4000 ;
        RECT  18.8650 0.7600 18.9850 1.5200 ;
        RECT  18.2050 1.2800 18.3250 2.1700 ;
        RECT  18.0850 0.5900 18.2050 0.8800 ;
        RECT  17.3650 1.2800 17.4850 2.1700 ;
        RECT  17.2450 0.5900 17.3650 0.8800 ;
        RECT  16.5250 1.2800 16.6450 2.1700 ;
        RECT  16.4050 0.5900 16.5250 1.4000 ;
        RECT  15.5650 0.7600 16.5250 0.8800 ;
        RECT  15.6850 1.2800 15.8050 2.1700 ;
        RECT  15.5650 0.5900 15.6850 0.8800 ;
        RECT  14.8450 1.2800 14.9650 2.1700 ;
        RECT  14.7250 0.5900 14.8450 0.8300 ;
        RECT  14.5450 0.7100 14.8450 0.8300 ;
        RECT  14.5450 0.7100 14.6650 1.4000 ;
        RECT  13.8850 0.7600 14.6650 0.8800 ;
        RECT  14.0050 1.2800 14.1250 2.1700 ;
        RECT  13.8850 0.5900 14.0050 0.8800 ;
        RECT  13.1650 1.2800 13.2850 2.1700 ;
        RECT  13.0450 0.5900 13.1650 0.8300 ;
        RECT  12.8650 0.7100 13.1650 0.8300 ;
        RECT  12.8650 0.7100 12.9850 1.4000 ;
        RECT  12.2050 0.7600 12.9850 0.8800 ;
        RECT  12.3250 1.2800 12.4450 2.1700 ;
        RECT  12.2050 0.5900 12.3250 0.8800 ;
        RECT  11.6700 0.8850 11.8200 1.1450 ;
        RECT  11.6650 0.9200 11.7900 1.4000 ;
        RECT  11.4850 1.5200 11.7850 1.6400 ;
        RECT  11.6650 0.9200 11.7850 1.6400 ;
        RECT  11.3650 0.9200 11.8200 1.0400 ;
        RECT  11.4850 1.5200 11.6050 2.1700 ;
        RECT  11.3650 0.5900 11.4850 1.0400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 19.7200 0.1800 ;
        RECT  19.3450 -0.1800 19.4650 0.6400 ;
        RECT  18.5050 -0.1800 18.6250 0.6400 ;
        RECT  17.6650 -0.1800 17.7850 0.6400 ;
        RECT  16.8250 -0.1800 16.9450 0.6400 ;
        RECT  15.9850 -0.1800 16.1050 0.6400 ;
        RECT  15.1450 -0.1800 15.2650 0.6400 ;
        RECT  14.3050 -0.1800 14.4250 0.6400 ;
        RECT  13.4650 -0.1800 13.5850 0.6400 ;
        RECT  12.6250 -0.1800 12.7450 0.6400 ;
        RECT  11.7850 -0.1800 11.9050 0.6400 ;
        RECT  10.8850 0.4600 11.1250 0.5800 ;
        RECT  10.8850 -0.1800 11.0050 0.5800 ;
        RECT  10.0450 0.4600 10.2850 0.5800 ;
        RECT  10.0450 -0.1800 10.1650 0.5800 ;
        RECT  9.2050 0.4600 9.4450 0.5800 ;
        RECT  9.2050 -0.1800 9.3250 0.5800 ;
        RECT  8.3650 0.4600 8.6050 0.5800 ;
        RECT  8.3650 -0.1800 8.4850 0.5800 ;
        RECT  7.5250 0.4600 7.7650 0.5800 ;
        RECT  7.5250 -0.1800 7.6450 0.5800 ;
        RECT  6.6850 0.4600 6.9250 0.5800 ;
        RECT  6.6850 -0.1800 6.8050 0.5800 ;
        RECT  5.9050 -0.1800 6.0250 0.6400 ;
        RECT  4.8250 -0.1800 4.9450 0.6650 ;
        RECT  3.3250 -0.1800 3.4450 0.6600 ;
        RECT  1.8450 -0.1800 1.9650 0.6600 ;
        RECT  0.3650 -0.1800 0.4850 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 19.7200 2.7900 ;
        RECT  19.4650 1.5200 19.5850 2.7900 ;
        RECT  18.6250 1.5200 18.7450 2.7900 ;
        RECT  17.7850 1.5200 17.9050 2.7900 ;
        RECT  16.9450 1.5200 17.0650 2.7900 ;
        RECT  16.1050 1.5200 16.2250 2.7900 ;
        RECT  15.2650 1.5200 15.3850 2.7900 ;
        RECT  14.4250 1.5200 14.5450 2.7900 ;
        RECT  13.5850 1.5200 13.7050 2.7900 ;
        RECT  12.7450 1.5200 12.8650 2.7900 ;
        RECT  11.9050 1.5200 12.0250 2.7900 ;
        RECT  11.0050 1.9000 11.2450 2.1100 ;
        RECT  11.0050 1.9000 11.1250 2.7900 ;
        RECT  9.1650 1.9000 9.4050 2.0200 ;
        RECT  9.1650 1.9000 9.2850 2.7900 ;
        RECT  7.5050 2.0550 7.7450 2.1750 ;
        RECT  7.5050 2.0550 7.6250 2.7900 ;
        RECT  6.1050 2.0100 6.3450 2.1300 ;
        RECT  6.1050 2.0100 6.2250 2.7900 ;
        RECT  5.2050 1.5100 5.3250 2.7900 ;
        RECT  4.3050 2.2300 4.4250 2.7900 ;
        RECT  3.5850 2.2300 3.7050 2.7900 ;
        RECT  2.7450 2.2300 2.8650 2.7900 ;
        RECT  1.9050 2.2300 2.0250 2.7900 ;
        RECT  1.0650 2.2300 1.1850 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.4450 1.4000 11.3650 1.4000 11.3650 1.7800 10.5700 1.7800 10.5700 2.2500
                 9.5250 2.2500 9.5250 1.7800 9.0450 1.7800 9.0450 2.2500 7.8650 2.2500 7.8650 1.9350
                 6.5400 1.9350 6.5400 1.8900 5.4450 1.8900 5.4450 1.3900 4.9050 1.3900 4.9050 1.9500
                 4.7850 1.9500 4.7850 1.6200 4.0650 1.6200 4.0650 1.9500 3.9450 1.9500 3.9450 1.6200
                 3.2250 1.6200 3.2250 1.9500 3.1050 1.9500 3.1050 1.6200 2.3850 1.6200 2.3850 1.9500
                 2.2650 1.9500 2.2650 1.6200 1.5450 1.6200 1.5450 1.9500 1.4250 1.9500 1.4250 1.6200
                 0.7050 1.6200 0.7050 1.9500 0.5850 1.9500 0.5850 1.4050 0.7050 1.4050 0.7050 1.5000
                 0.9450 1.5000 0.9450 0.6000 1.1850 0.6000 1.1850 0.7200 1.0650 0.7200 1.0650 1.5000
                 1.4250 1.5000 1.4250 1.4800 1.5450 1.4800 1.5450 1.5000 2.2650 1.5000 2.2650 1.4800
                 2.3850 1.4800 2.3850 1.5000 2.6050 1.5000 2.6050 0.7200 2.5850 0.7200 2.5850 0.6000
                 2.8250 0.6000 2.8250 0.7200 2.7250 0.7200 2.7250 1.5000 3.9450 1.5000 3.9450 1.4600
                 4.0650 1.4600 4.0650 1.5000 4.3450 1.5000 4.3450 0.7200 4.1250 0.7200 4.1250 0.6000
                 4.4650 0.6000 4.4650 1.5000 4.7850 1.5000 4.7850 1.2700 5.5650 1.2700 5.5650 1.7700
                 6.6600 1.7700 6.6600 1.8150 7.9850 1.8150 7.9850 2.1300 8.9250 2.1300 8.9250 1.6600
                 9.6450 1.6600 9.6450 2.1300 10.4500 2.1300 10.4500 1.6600 11.2450 1.6600
                 11.2450 1.2800 11.3250 1.2800 11.3250 1.1600 11.4450 1.1600 ;
        POLYGON  11.1250 1.1700 11.1050 1.1700 11.1050 1.5400 10.2250 1.5400 10.2250 2.0100
                 10.1050 2.0100 10.1050 1.5400 8.5450 1.5400 8.5450 2.0100 8.4250 2.0100 8.4250 1.5400
                 7.0450 1.5400 7.0450 1.6950 6.8050 1.6950 6.8050 1.5750 6.9250 1.5750 6.9250 1.4200
                 10.9850 1.4200 10.9850 0.8200 6.3250 0.8200 6.3250 0.5200 6.4450 0.5200 6.4450 0.7000
                 7.1650 0.7000 7.1650 0.5200 7.2850 0.5200 7.2850 0.7000 8.0050 0.7000 8.0050 0.5200
                 8.1250 0.5200 8.1250 0.7000 8.8450 0.7000 8.8450 0.5200 8.9650 0.5200 8.9650 0.7000
                 9.6850 0.7000 9.6850 0.5150 9.8050 0.5150 9.8050 0.7000 10.5250 0.7000 10.5250 0.5150
                 10.6450 0.5150 10.6450 0.7000 11.1050 0.7000 11.1050 0.9300 11.1250 0.9300 ;
        POLYGON  10.0050 1.3000 5.8050 1.3000 5.8050 1.6500 5.6850 1.6500 5.6850 1.1200 5.3050 1.1200
                 5.3050 0.6500 5.5450 0.6500 5.5450 1.0000 5.8050 1.0000 5.8050 1.1800 10.0050 1.1800 ;
        POLYGON  2.4850 1.3600 1.2850 1.3600 1.2850 1.0850 1.4050 1.0850 1.4050 1.2400 2.3650 1.2400
                 2.3650 1.0900 2.4850 1.0900 ;
    END
END TBUFX20

MACRO TBUFX2
    CLASS CORE ;
    FOREIGN TBUFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9450 0.7800 1.1850 0.9000 ;
        RECT  0.4450 0.8600 1.0650 0.9800 ;
        RECT  0.4450 0.8600 0.5650 1.2200 ;
        RECT  0.3050 0.9400 0.5650 1.0900 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1750 0.9800 2.4150 1.1000 ;
        RECT  1.1150 1.7600 2.2950 1.8800 ;
        RECT  2.1750 0.9800 2.2950 1.8800 ;
        RECT  0.8850 1.6700 1.2350 1.7900 ;
        RECT  0.8850 1.5200 1.1450 1.7900 ;
        RECT  0.8850 1.1000 1.0050 1.7900 ;
        RECT  0.7250 1.1000 1.0050 1.2200 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0950 1.1450 3.2150 1.8800 ;
        RECT  2.9700 0.8850 3.1200 1.2650 ;
        RECT  2.9350 0.5900 3.0550 1.0250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.3550 -0.1800 3.4750 0.6400 ;
        RECT  2.4550 0.5000 2.6950 0.6200 ;
        RECT  2.4550 -0.1800 2.5750 0.6200 ;
        RECT  1.6750 -0.1800 1.7950 0.6800 ;
        RECT  0.8650 -0.1800 0.9850 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.5150 1.3400 3.6350 2.7900 ;
        RECT  2.5550 2.2400 2.7950 2.7900 ;
        RECT  0.9450 2.2400 1.1850 2.7900 ;
        RECT  0.1350 1.5800 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1550 2.2500 2.9150 2.2500 2.9150 2.1200 0.5550 2.1200 0.5550 1.4600 0.0650 1.4600
                 0.0650 0.6200 0.2250 0.6200 0.2250 0.4000 0.3450 0.4000 0.3450 0.7400 0.1850 0.7400
                 0.1850 1.3400 0.6750 1.3400 0.6750 2.0000 3.0350 2.0000 3.0350 2.1300 3.1550 2.1300 ;
        POLYGON  2.7150 1.1500 2.5950 1.1500 2.5950 0.8600 2.0550 0.8600 2.0550 1.6400 1.8150 1.6400
                 1.8150 1.5200 1.9350 1.5200 1.9350 0.7400 2.0950 0.7400 2.0950 0.4400 2.2150 0.4400
                 2.2150 0.7400 2.7150 0.7400 ;
        POLYGON  1.8150 1.0200 1.5450 1.0200 1.5450 1.5200 1.6650 1.5200 1.6650 1.6400 1.4250 1.6400
                 1.4250 0.6600 1.2850 0.6600 1.2850 0.4000 1.4050 0.4000 1.4050 0.5400 1.5450 0.5400
                 1.5450 0.9000 1.8150 0.9000 ;
    END
END TBUFX2

MACRO TBUFX16
    CLASS CORE ;
    FOREIGN TBUFX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 16.5300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.2184  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.5400  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.4044  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5150 0.8500 1.6350 1.1000 ;
        RECT  0.5550 0.8500 1.6350 0.9700 ;
        RECT  0.3600 0.8850 0.6750 1.1250 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8550 1.1850 9.0950 1.3050 ;
        RECT  8.8550 1.0000 8.9750 1.3050 ;
        RECT  5.5150 1.0000 8.9750 1.1200 ;
        RECT  5.5150 0.7600 5.6350 1.1200 ;
        RECT  4.9350 0.7600 5.6350 0.8800 ;
        RECT  4.9350 0.4100 5.0550 0.8800 ;
        RECT  4.3350 0.4100 5.0550 0.5300 ;
        RECT  3.8550 0.7950 4.4550 0.9150 ;
        RECT  4.3350 0.4100 4.4550 0.9150 ;
        RECT  4.1200 0.7950 4.2400 1.1500 ;
        RECT  3.8550 0.3600 3.9750 0.9150 ;
        RECT  3.1550 0.3600 3.9750 0.4800 ;
        RECT  2.4500 0.7100 3.2750 0.8300 ;
        RECT  3.1550 0.3600 3.2750 0.8300 ;
        RECT  2.7150 0.7100 2.8350 1.1200 ;
        RECT  2.4500 0.3600 2.5700 0.8300 ;
        RECT  1.7550 0.3600 2.5700 0.4800 ;
        RECT  1.7550 0.9400 2.0150 1.0900 ;
        RECT  1.1750 1.2200 1.8750 1.3400 ;
        RECT  1.7550 0.3600 1.8750 1.3400 ;
        RECT  0.7950 1.1500 1.2950 1.2700 ;
        RECT  1.1750 1.0900 1.2950 1.3400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  15.6950 1.3200 15.8150 2.2100 ;
        RECT  15.6750 0.5900 15.7950 1.4400 ;
        RECT  9.9300 1.3200 15.8150 1.4400 ;
        RECT  13.9950 0.7600 15.7950 0.8800 ;
        RECT  14.8550 1.3200 14.9750 2.2100 ;
        RECT  14.8350 0.5900 14.9550 0.8800 ;
        RECT  14.0150 1.3200 14.1350 2.2100 ;
        RECT  13.9950 0.5900 14.1150 0.8800 ;
        RECT  13.1750 1.3200 13.2950 2.2100 ;
        RECT  13.1550 0.5900 13.2750 1.4400 ;
        RECT  12.3150 0.7600 13.2750 0.8800 ;
        RECT  12.3350 1.3200 12.4550 2.2100 ;
        RECT  12.3150 0.5900 12.4350 0.8800 ;
        RECT  11.4950 1.3200 11.6150 2.2100 ;
        RECT  11.4750 0.5900 11.5950 0.8300 ;
        RECT  11.2950 0.7100 11.5950 0.8300 ;
        RECT  11.2950 0.7100 11.4150 1.4400 ;
        RECT  10.6350 0.7600 11.4150 0.8800 ;
        RECT  10.6550 1.3200 10.7750 2.2100 ;
        RECT  10.6350 0.5900 10.7550 0.8800 ;
        RECT  9.9300 1.1750 10.0800 1.4400 ;
        RECT  9.9300 0.9600 10.0500 1.6800 ;
        RECT  9.8150 1.5600 9.9350 2.2100 ;
        RECT  9.7950 0.9600 10.0500 1.0800 ;
        RECT  9.7950 0.5900 9.9150 1.0800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 16.5300 0.1800 ;
        RECT  16.0950 -0.1800 16.2150 0.6400 ;
        RECT  15.2550 -0.1800 15.3750 0.6400 ;
        RECT  14.4150 -0.1800 14.5350 0.6400 ;
        RECT  13.5750 -0.1800 13.6950 0.6400 ;
        RECT  12.7350 -0.1800 12.8550 0.6400 ;
        RECT  11.8950 -0.1800 12.0150 0.6400 ;
        RECT  11.0550 -0.1800 11.1750 0.6400 ;
        RECT  10.2150 -0.1800 10.3350 0.6400 ;
        RECT  9.3750 -0.1800 9.4950 0.6400 ;
        RECT  8.5350 -0.1800 8.6550 0.6400 ;
        RECT  7.6950 -0.1800 7.8150 0.6400 ;
        RECT  6.8550 -0.1800 6.9750 0.6400 ;
        RECT  6.0150 -0.1800 6.1350 0.6400 ;
        RECT  5.1750 -0.1800 5.2950 0.6400 ;
        RECT  4.0950 -0.1800 4.2150 0.6750 ;
        RECT  2.6950 0.4700 2.9350 0.5900 ;
        RECT  2.6950 -0.1800 2.8150 0.5900 ;
        RECT  0.9550 -0.1800 1.0750 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 16.5300 2.7900 ;
        RECT  16.1150 1.5600 16.2350 2.7900 ;
        RECT  15.2750 1.5600 15.3950 2.7900 ;
        RECT  14.4350 1.5600 14.5550 2.7900 ;
        RECT  13.5950 1.5600 13.7150 2.7900 ;
        RECT  12.7550 1.5600 12.8750 2.7900 ;
        RECT  11.9150 1.5600 12.0350 2.7900 ;
        RECT  11.0750 1.5600 11.1950 2.7900 ;
        RECT  10.2350 1.5600 10.3550 2.7900 ;
        RECT  8.9950 1.9600 9.2350 2.0800 ;
        RECT  8.9950 1.9600 9.1150 2.7900 ;
        RECT  7.7150 1.9600 7.9550 2.0800 ;
        RECT  7.7150 1.9600 7.8350 2.7900 ;
        RECT  6.4350 1.9600 6.6750 2.0800 ;
        RECT  6.4350 1.9600 6.5550 2.7900 ;
        RECT  4.7350 1.5300 4.8550 2.7900 ;
        RECT  4.6150 1.5300 4.8550 1.9300 ;
        RECT  3.8350 1.7200 3.9550 2.7900 ;
        RECT  2.9350 2.2300 3.0550 2.7900 ;
        RECT  2.0350 1.7200 2.1550 2.7900 ;
        RECT  1.1350 2.2300 1.2550 2.7900 ;
        RECT  0.2350 1.7200 0.3550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.7950 1.4400 9.6950 1.4400 9.6950 1.8400 8.7750 1.8400 8.7750 2.2500 8.0750 2.2500
                 8.0750 1.8400 7.5450 1.8400 7.5450 2.2500 6.8950 2.2500 6.8950 1.8400 6.2750 1.8400
                 6.2750 2.2500 4.9750 2.2500 4.9750 1.4100 4.3750 1.4100 4.3750 1.9900 4.2550 1.9900
                 4.2550 1.6000 3.5350 1.6000 3.5350 1.9500 3.4150 1.9500 3.4150 1.6000 2.5750 1.6000
                 2.5750 1.9800 2.4550 1.9800 2.4550 1.6000 1.7350 1.6000 1.7350 1.9500 1.6150 1.9500
                 1.6150 1.6000 0.7750 1.6000 0.7750 2.2100 0.6550 2.2100 0.6550 1.6000 0.1200 1.6000
                 0.1200 0.6450 0.3150 0.6450 0.3150 0.5250 0.4350 0.5250 0.4350 0.7650 0.2400 0.7650
                 0.2400 1.4800 1.6150 1.4800 1.6150 1.4600 1.7350 1.4600 1.7350 1.4800 2.1350 1.4800
                 2.1350 0.7200 1.9950 0.7200 1.9950 0.6000 2.2550 0.6000 2.2550 1.4800 3.6150 1.4800
                 3.6150 0.7200 3.3950 0.7200 3.3950 0.6000 3.7350 0.6000 3.7350 1.4800 4.2550 1.4800
                 4.2550 1.2900 5.0950 1.2900 5.0950 2.1300 6.1550 2.1300 6.1550 1.7200 7.0150 1.7200
                 7.0150 2.1300 7.4250 2.1300 7.4250 1.7200 8.1950 1.7200 8.1950 2.1300 8.6550 2.1300
                 8.6550 1.7200 9.5750 1.7200 9.5750 1.3200 9.6750 1.3200 9.6750 1.2000 9.7950 1.2000 ;
        POLYGON  9.4550 1.2250 9.3350 1.2250 9.3350 1.6000 8.5350 1.6000 8.5350 2.0100 8.4150 2.0100
                 8.4150 1.6000 7.2550 1.6000 7.2550 2.0100 7.1350 2.0100 7.1350 1.6000 6.0350 1.6000
                 6.0350 2.0100 5.7950 2.0100 5.7950 1.6800 5.9150 1.6800 5.9150 1.4800 9.2150 1.4800
                 9.2150 0.8800 5.7550 0.8800 5.7550 0.6400 5.5950 0.6400 5.5950 0.4000 5.7150 0.4000
                 5.7150 0.5200 5.8750 0.5200 5.8750 0.7600 6.4350 0.7600 6.4350 0.5050 6.5550 0.5050
                 6.5550 0.7600 7.2750 0.7600 7.2750 0.5050 7.3950 0.5050 7.3950 0.7600 8.1150 0.7600
                 8.1150 0.5050 8.2350 0.5050 8.2350 0.7600 8.9550 0.7600 8.9550 0.5050 9.0750 0.5050
                 9.0750 0.7600 9.3350 0.7600 9.3350 1.1050 9.4550 1.1050 ;
        POLYGON  8.4550 1.3600 5.5150 1.3600 5.5150 1.9300 5.2750 1.9300 5.2750 1.1200 4.5750 1.1200
                 4.5750 0.6500 4.8150 0.6500 4.8150 1.0000 5.3950 1.0000 5.3950 1.2400 8.4550 1.2400 ;
        POLYGON  3.4950 1.3600 2.3750 1.3600 2.3750 1.1200 2.4950 1.1200 2.4950 1.2400 3.2550 1.2400
                 3.2550 0.9500 3.4950 0.9500 ;
    END
END TBUFX16

MACRO TBUFX12
    CLASS CORE ;
    FOREIGN TBUFX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.4700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.1584  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.3667  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 0.8650 1.3350 1.1050 ;
        RECT  0.5350 0.9700 1.3350 1.0900 ;
        RECT  0.5950 0.9400 0.8550 1.0900 ;
        RECT  0.5350 0.9700 0.6550 1.2300 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0200 1.1800 6.9950 1.3000 ;
        RECT  6.8750 1.0600 6.9950 1.3000 ;
        RECT  4.0200 1.0200 4.1750 1.3000 ;
        RECT  3.4950 0.9000 4.1400 1.0200 ;
        RECT  3.9350 1.0200 4.1750 1.1400 ;
        RECT  3.4950 0.3600 3.6150 1.0200 ;
        RECT  2.7950 0.3600 3.6150 0.4800 ;
        RECT  2.1550 0.7600 2.9150 0.8800 ;
        RECT  2.7950 0.3600 2.9150 0.8800 ;
        RECT  2.2350 0.7600 2.4750 1.0450 ;
        RECT  2.1550 0.3650 2.2750 0.8800 ;
        RECT  1.4550 0.3650 2.2750 0.4850 ;
        RECT  0.9150 1.2250 1.5750 1.3450 ;
        RECT  1.4550 0.3650 1.5750 1.3450 ;
        RECT  1.1750 1.2250 1.4350 1.3800 ;
        RECT  0.7950 1.2100 1.0350 1.3300 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.7950 1.4400 11.9150 2.2100 ;
        RECT  11.7750 0.5900 11.8950 0.8300 ;
        RECT  11.6150 1.4400 11.9150 1.5600 ;
        RECT  11.5950 0.7100 11.8950 0.8300 ;
        RECT  7.7550 1.3200 11.7350 1.4400 ;
        RECT  11.5950 0.7100 11.7150 1.4400 ;
        RECT  10.0950 0.7600 11.7150 0.8800 ;
        RECT  10.9550 1.3200 11.0750 2.2100 ;
        RECT  10.9350 0.5900 11.0550 0.8800 ;
        RECT  10.1150 1.3200 10.2350 2.2100 ;
        RECT  10.0950 0.5900 10.2150 0.8800 ;
        RECT  9.2750 1.3200 9.3950 2.2100 ;
        RECT  9.2550 0.5900 9.3750 0.8300 ;
        RECT  9.0750 0.7100 9.3750 0.8300 ;
        RECT  9.0750 0.7100 9.1950 1.4400 ;
        RECT  8.4150 0.7600 9.1950 0.8800 ;
        RECT  8.4350 1.3200 8.5550 2.2100 ;
        RECT  8.4150 0.5900 8.5350 0.8800 ;
        RECT  7.7550 1.1750 8.0500 1.4400 ;
        RECT  7.5950 1.5400 7.8750 1.6600 ;
        RECT  7.7550 0.7100 7.8750 1.6600 ;
        RECT  7.5750 0.7100 7.8750 0.8300 ;
        RECT  7.5950 1.5400 7.7150 2.2100 ;
        RECT  7.5750 0.5900 7.6950 0.8300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.4700 0.1800 ;
        RECT  12.1950 -0.1800 12.3150 0.6400 ;
        RECT  11.3550 -0.1800 11.4750 0.6400 ;
        RECT  10.5150 -0.1800 10.6350 0.6400 ;
        RECT  9.6750 -0.1800 9.7950 0.6400 ;
        RECT  8.8350 -0.1800 8.9550 0.6400 ;
        RECT  7.9950 -0.1800 8.1150 0.6400 ;
        RECT  7.1550 -0.1800 7.2750 0.6400 ;
        RECT  6.2550 0.4600 6.4950 0.5800 ;
        RECT  6.2550 -0.1800 6.3750 0.5800 ;
        RECT  5.4150 0.4600 5.6550 0.5800 ;
        RECT  5.4150 -0.1800 5.5350 0.5800 ;
        RECT  4.5750 0.4600 4.8150 0.5800 ;
        RECT  4.5750 -0.1800 4.6950 0.5800 ;
        RECT  3.7350 0.5200 3.9750 0.6400 ;
        RECT  3.8550 -0.1800 3.9750 0.6400 ;
        RECT  2.3950 0.5200 2.6350 0.6400 ;
        RECT  2.5150 -0.1800 2.6350 0.6400 ;
        RECT  0.7150 -0.1800 0.8350 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.4700 2.7900 ;
        RECT  12.2150 1.5600 12.3350 2.7900 ;
        RECT  11.3750 1.5600 11.4950 2.7900 ;
        RECT  10.5350 1.5600 10.6550 2.7900 ;
        RECT  9.6950 1.5600 9.8150 2.7900 ;
        RECT  8.8550 1.5600 8.9750 2.7900 ;
        RECT  8.0150 1.5600 8.1350 2.7900 ;
        RECT  7.1750 1.9000 7.2950 2.7900 ;
        RECT  5.6550 2.0150 5.8950 2.1350 ;
        RECT  5.6550 2.0150 5.7750 2.7900 ;
        RECT  4.2350 2.2250 4.3550 2.7900 ;
        RECT  3.3550 2.2250 3.4750 2.7900 ;
        RECT  2.5150 2.2250 2.6350 2.7900 ;
        RECT  1.5750 2.2300 1.6950 2.7900 ;
        RECT  0.5550 2.0300 0.7950 2.1500 ;
        RECT  0.5550 2.0300 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.5950 1.4200 7.4750 1.4200 7.4750 1.7800 6.7750 1.7800 6.7750 2.2050 6.0400 2.2050
                 6.0400 1.8950 4.7150 1.8950 4.7150 1.8650 3.8350 1.8650 3.8350 1.6200 3.0550 1.6200
                 3.0550 1.6400 2.8150 1.6400 2.8150 1.6200 2.2150 1.6200 2.2150 1.6400 1.9750 1.6400
                 1.9750 1.6200 1.2750 1.6200 1.2750 1.6700 1.0350 1.6700 1.0350 1.5500 1.1550 1.5500
                 1.1550 1.5000 1.6950 1.5000 1.6950 0.6050 1.9350 0.6050 1.9350 0.7250 1.8150 0.7250
                 1.8150 1.5000 3.2550 1.5000 3.2550 0.7200 3.0350 0.7200 3.0350 0.6000 3.3750 0.6000
                 3.3750 1.5000 3.9550 1.5000 3.9550 1.7450 4.8350 1.7450 4.8350 1.7750 6.1600 1.7750
                 6.1600 2.0850 6.6550 2.0850 6.6550 1.6600 7.3550 1.6600 7.3550 1.3000 7.5950 1.3000 ;
        POLYGON  7.4150 1.1500 7.2350 1.1500 7.2350 1.5400 6.5350 1.5400 6.5350 1.9650 6.4150 1.9650
                 6.4150 1.5400 5.1950 1.5400 5.1950 1.6550 4.9550 1.6550 4.9550 1.5350 5.0750 1.5350
                 5.0750 1.4200 7.1150 1.4200 7.1150 0.9400 6.7350 0.9400 6.7350 0.8200 4.2600 0.8200
                 4.2600 0.7250 4.2150 0.7250 4.2150 0.4850 4.3350 0.4850 4.3350 0.6050 4.3800 0.6050
                 4.3800 0.7000 5.0550 0.7000 5.0550 0.4850 5.1750 0.4850 5.1750 0.7000 5.8950 0.7000
                 5.8950 0.4800 6.0150 0.4800 6.0150 0.7000 6.6900 0.7000 6.6900 0.6000 6.7350 0.6000
                 6.7350 0.4800 6.8550 0.4800 6.8550 0.8200 7.4150 0.8200 ;
        RECT  4.7950 0.9400 6.4350 1.0600 ;
        POLYGON  5.0350 2.2450 4.4750 2.2450 4.4750 2.1050 1.5600 2.1050 1.5600 1.9100 0.2550 1.9100
                 0.2550 2.1400 0.1350 2.1400 0.1350 1.4900 0.2950 1.4900 0.2950 0.6500 0.4150 0.6500
                 0.4150 1.6100 0.2550 1.6100 0.2550 1.7900 1.6800 1.7900 1.6800 1.9850 4.5950 1.9850
                 4.5950 2.1250 5.0350 2.1250 ;
        POLYGON  3.1350 1.2850 2.0550 1.2850 2.0550 1.3800 1.9350 1.3800 1.9350 1.1400 2.0550 1.1400
                 2.0550 1.1650 3.1350 1.1650 ;
    END
END TBUFX12

MACRO TBUFX1
    CLASS CORE ;
    FOREIGN TBUFX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3000 1.1600 1.2800 1.2800 ;
        RECT  0.6500 0.8850 0.8000 1.2800 ;
        RECT  0.3000 1.1600 0.4200 1.4000 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0150 0.3600 2.5150 0.4800 ;
        RECT  1.0800 0.4400 2.1350 0.5600 ;
        RECT  0.7000 1.4000 1.5200 1.5200 ;
        RECT  1.4000 0.9200 1.5200 1.5200 ;
        RECT  1.1750 1.4000 1.4350 1.6700 ;
        RECT  1.0800 0.9200 1.5200 1.0400 ;
        RECT  1.0800 0.4400 1.2000 1.0400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2650 0.7600 3.3850 1.6800 ;
        RECT  3.2250 1.5600 3.3450 2.2100 ;
        RECT  3.0550 0.7600 3.3850 0.8800 ;
        RECT  2.9150 0.6500 3.2150 0.8000 ;
        RECT  3.0950 0.6400 3.2150 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.6750 -0.1800 2.7950 0.6900 ;
        RECT  1.6550 -0.1800 1.8950 0.3200 ;
        RECT  0.8400 -0.1800 0.9600 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.8050 1.7000 2.9250 2.7900 ;
        RECT  0.9750 2.2700 1.2150 2.7900 ;
        RECT  0.1350 1.8500 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1450 1.4400 3.1050 1.4400 3.1050 1.5800 2.5950 1.5800 2.5950 2.1500 0.5550 2.1500
                 0.5550 1.8500 0.4600 1.8500 0.4600 1.6400 0.0600 1.6400 0.0600 0.9200 0.1400 0.9200
                 0.1400 0.6200 0.2600 0.6200 0.2600 1.0400 0.1800 1.0400 0.1800 1.5200 0.5800 1.5200
                 0.5800 1.7300 0.6750 1.7300 0.6750 2.0300 2.4750 2.0300 2.4750 1.4600 2.9850 1.4600
                 2.9850 1.2000 3.1450 1.2000 ;
        POLYGON  2.8650 1.3400 2.3550 1.3400 2.3550 1.6200 2.1450 1.6200 2.1450 1.7400 1.9050 1.7400
                 1.9050 1.6200 2.0250 1.6200 2.0250 1.5000 2.2350 1.5000 2.2350 0.8000 2.1350 0.8000
                 2.1350 0.6800 2.3750 0.6800 2.3750 0.8000 2.3550 0.8000 2.3550 1.2200 2.8650 1.2200 ;
        POLYGON  2.1150 1.3200 1.7600 1.3200 1.7600 1.9100 1.4550 1.9100 1.4550 1.7900 1.6400 1.7900
                 1.6400 0.8000 1.3200 0.8000 1.3200 0.6800 1.7600 0.6800 1.7600 1.2000 2.1150 1.2000 ;
    END
END TBUFX1

MACRO SMDFFHQX8
    CLASS CORE ;
    FOREIGN SMDFFHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.2100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 1.4450 2.7750 2.1900 ;
        RECT  2.6550 0.6650 2.7750 0.9050 ;
        RECT  2.6350 0.7850 2.7550 1.5650 ;
        RECT  0.0700 0.9050 2.7550 1.0250 ;
        RECT  1.8150 0.6650 1.9350 2.1900 ;
        RECT  0.9750 0.6650 1.0950 2.1850 ;
        RECT  0.1350 0.6650 0.2550 2.1850 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 1.1750 5.2050 1.3800 ;
        RECT  5.0850 1.0300 5.2050 1.3800 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6700 1.1600 9.9150 1.2800 ;
        RECT  9.6700 0.8850 9.7900 1.2800 ;
        RECT  9.6400 0.8850 9.7900 1.1450 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.3800 0.8850 11.5300 1.1450 ;
        RECT  11.2950 1.0250 11.4150 1.3850 ;
        END
    END SE
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.5950 1.2650 11.8350 1.3850 ;
        RECT  11.6700 0.8850 11.8200 1.1450 ;
        RECT  11.6700 0.8850 11.7900 1.3850 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.0500 1.2100 13.3550 1.4200 ;
        RECT  13.0500 1.2100 13.3250 1.4450 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.4950 0.9700 13.6150 1.2100 ;
        RECT  12.5350 0.9700 13.6150 1.0900 ;
        RECT  12.7750 0.9400 13.0350 1.0900 ;
        RECT  12.3150 1.0000 12.6550 1.1200 ;
        RECT  12.1950 1.2650 12.4350 1.3850 ;
        RECT  12.3150 1.0000 12.4350 1.3850 ;
        END
    END S0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.2100 0.1800 ;
        RECT  13.3350 -0.1800 13.4550 0.8200 ;
        RECT  12.0550 -0.1800 12.1750 0.6400 ;
        RECT  9.8550 -0.1800 9.9750 0.7650 ;
        RECT  7.5850 0.4100 7.8250 0.5300 ;
        RECT  7.7050 -0.1800 7.8250 0.5300 ;
        RECT  5.3250 0.3100 5.5650 0.4300 ;
        RECT  5.4450 -0.1800 5.5650 0.4300 ;
        RECT  3.9150 -0.1800 4.0350 0.6500 ;
        RECT  3.0750 -0.1800 3.1950 0.6500 ;
        RECT  2.2350 -0.1800 2.3550 0.6550 ;
        RECT  1.3950 -0.1800 1.5150 0.6550 ;
        RECT  0.5550 -0.1800 0.6750 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.2100 2.7900 ;
        RECT  13.1350 1.8050 13.2550 2.7900 ;
        RECT  11.7550 1.7450 11.8750 2.7900 ;
        RECT  9.7950 1.7500 9.9150 2.7900 ;
        RECT  7.5850 2.0100 7.8250 2.1300 ;
        RECT  7.5850 2.0100 7.7050 2.7900 ;
        RECT  5.6850 1.9800 5.8050 2.7900 ;
        RECT  3.9150 1.5400 4.0350 2.7900 ;
        RECT  3.0750 1.5400 3.1950 2.7900 ;
        RECT  2.2350 1.4450 2.3550 2.7900 ;
        RECT  1.3950 1.4450 1.5150 2.7900 ;
        RECT  0.5550 1.4450 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.8750 0.8200 13.8550 0.8200 13.8550 1.6850 13.7750 1.6850 13.7750 1.8050
                 13.6550 1.8050 13.6550 1.6850 12.6350 1.6850 12.6350 1.2400 12.7550 1.2400
                 12.7550 1.5650 13.7350 1.5650 13.7350 0.7000 13.7550 0.7000 13.7550 0.5800
                 13.8750 0.5800 ;
        POLYGON  12.8150 0.8200 12.4150 0.8200 12.4150 0.8800 12.0750 0.8800 12.0750 1.5050
                 12.5150 1.5050 12.5150 2.2100 12.3950 2.2100 12.3950 1.6250 11.0350 1.6250
                 11.0350 1.8200 10.9150 1.8200 10.9150 1.4900 11.0550 1.4900 11.0550 0.7650
                 11.0350 0.7650 11.0350 0.6450 11.2750 0.6450 11.2750 0.7650 11.1750 0.7650
                 11.1750 1.5050 11.9550 1.5050 11.9550 0.7600 12.2950 0.7600 12.2950 0.7000
                 12.6950 0.7000 12.6950 0.5600 12.8150 0.5600 ;
        POLYGON  11.7150 0.7650 11.4750 0.7650 11.4750 0.5250 10.9150 0.5250 10.9150 0.8850
                 10.9350 0.8850 10.9350 1.3700 10.7950 1.3700 10.7950 1.9700 11.3950 1.9700
                 11.3950 2.2100 11.2750 2.2100 11.2750 2.0900 10.6750 2.0900 10.6750 1.2700
                 10.3950 1.2700 10.3950 1.3900 10.2750 1.3900 10.2750 1.1500 10.8150 1.1500
                 10.8150 1.0050 10.7950 1.0050 10.7950 0.4050 11.5950 0.4050 11.5950 0.6450
                 11.7150 0.6450 ;
        POLYGON  10.6750 0.7700 10.5550 0.7700 10.5550 1.0050 10.1550 1.0050 10.1550 1.5100
                 10.5550 1.5100 10.5550 2.1400 10.4350 2.1400 10.4350 1.6300 9.1050 1.6300
                 9.1050 1.9300 8.9850 1.9300 8.9850 1.4400 9.0250 1.4400 9.0250 0.7200 8.9850 0.7200
                 8.9850 0.6000 9.2250 0.6000 9.2250 0.7200 9.1450 0.7200 9.1450 1.5100 10.0350 1.5100
                 10.0350 0.8850 10.4350 0.8850 10.4350 0.6500 10.6750 0.6500 ;
        POLYGON  9.5550 0.7650 9.4350 0.7650 9.4350 0.4800 8.8650 0.4800 8.8650 1.0800 8.9050 1.0800
                 8.9050 1.3200 8.8650 1.3200 8.8650 2.0500 9.3150 2.0500 9.3150 1.9300 9.5550 1.9300
                 9.5550 2.0500 9.4350 2.0500 9.4350 2.1700 8.7450 2.1700 8.7450 0.4800 8.2650 0.4800
                 8.2650 0.9200 8.3850 0.9200 8.3850 1.0400 8.1450 1.0400 8.1450 0.7700 7.3450 0.7700
                 7.3450 0.4800 6.8650 0.4800 6.8650 0.8400 6.9850 0.8400 6.9850 1.1200 6.8650 1.1200
                 6.8650 0.9600 6.7450 0.9600 6.7450 0.3600 7.4650 0.3600 7.4650 0.6500 8.1450 0.6500
                 8.1450 0.3600 9.5550 0.3600 ;
        POLYGON  8.6250 1.9300 8.5050 1.9300 8.5050 1.2800 7.4850 1.2800 7.4850 1.2500 7.3650 1.2500
                 7.3650 1.1300 7.6050 1.1300 7.6050 1.1600 8.5050 1.1600 8.5050 0.7200 8.3850 0.7200
                 8.3850 0.6000 8.6250 0.6000 ;
        POLYGON  8.3450 2.2500 8.2250 2.2500 8.2250 1.8900 7.2850 1.8900 7.2850 2.1700 5.9450 2.1700
                 5.9450 0.9100 4.8250 0.9100 4.8250 1.5000 5.3050 1.5000 5.3050 1.6200 4.7050 1.6200
                 4.7050 0.6000 4.9650 0.6000 4.9650 0.7900 6.0650 0.7900 6.0650 2.0500 6.6250 2.0500
                 6.6250 1.3200 6.5250 1.3200 6.5250 1.0800 6.6450 1.0800 6.6450 1.2000 6.7450 1.2000
                 6.7450 2.0500 7.1650 2.0500 7.1650 1.7700 8.3450 1.7700 ;
        POLYGON  8.0250 1.0400 7.7250 1.0400 7.7250 1.0100 7.2250 1.0100 7.2250 1.6500 7.1050 1.6500
                 7.1050 0.7200 6.9850 0.7200 6.9850 0.6000 7.2250 0.6000 7.2250 0.8900 7.8450 0.8900
                 7.8450 0.9200 8.0250 0.9200 ;
        POLYGON  6.5050 1.9300 6.3850 1.9300 6.3850 1.5600 6.2850 1.5600 6.2850 0.6700 5.0850 0.6700
                 5.0850 0.4800 4.2750 0.4800 4.2750 1.1800 4.1550 1.1800 4.1550 0.3600 5.2050 0.3600
                 5.2050 0.5500 6.2850 0.5500 6.2850 0.5400 6.4050 0.5400 6.4050 1.4400 6.5050 1.4400 ;
        POLYGON  5.7250 1.8600 4.4550 1.8600 4.4550 2.1900 4.3350 2.1900 4.3350 1.5400 4.3950 1.5400
                 4.3950 1.4200 3.6150 1.4200 3.6150 2.1900 3.4950 2.1900 3.4950 1.2250 2.8750 1.2250
                 2.8750 1.1050 3.4950 1.1050 3.4950 0.6000 3.6150 0.6000 3.6150 1.3000 4.3950 1.3000
                 4.3950 0.6000 4.5150 0.6000 4.5150 1.7400 5.6050 1.7400 5.6050 1.0700 5.7250 1.0700 ;
    END
END SMDFFHQX8

MACRO SMDFFHQX4
    CLASS CORE ;
    FOREIGN SMDFFHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8350 1.5300 2.2350 1.6500 ;
        RECT  1.8550 0.6600 1.9750 0.9000 ;
        RECT  1.8350 0.7800 1.9550 1.6500 ;
        RECT  0.9400 1.3150 1.9550 1.4350 ;
        RECT  1.0350 1.3150 1.2750 1.6500 ;
        RECT  0.9400 1.1750 1.1550 1.4350 ;
        RECT  1.0350 0.7800 1.1550 1.6500 ;
        RECT  1.0150 0.6600 1.1350 0.9000 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0200 0.5100 1.4700 ;
        RECT  0.3750 0.9150 0.4950 1.4700 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3200 1.0600 7.5250 1.4400 ;
        RECT  7.4050 1.0500 7.5250 1.4400 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0600 0.8000 9.2100 1.2000 ;
        RECT  9.0400 0.8250 9.1600 1.2400 ;
        END
    END SE
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3800 0.7600 9.5000 1.2400 ;
        RECT  9.3500 0.7600 9.5000 1.2150 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.2100 10.9400 1.3450 ;
        RECT  10.4550 1.2100 10.7150 1.3800 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0800 0.9700 11.2000 1.2100 ;
        RECT  9.9750 0.9700 11.2000 1.0900 ;
        RECT  10.7450 0.9400 11.0050 1.0900 ;
        RECT  9.9750 0.9700 10.0950 1.3200 ;
        RECT  9.8600 1.2000 9.9800 1.4400 ;
        END
    END S0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  10.9200 -0.1800 11.0400 0.8200 ;
        RECT  9.4950 -0.1800 9.6150 0.6400 ;
        RECT  7.5050 -0.1800 7.6250 0.8100 ;
        RECT  5.2750 -0.1800 5.5150 0.3700 ;
        RECT  3.1150 0.4300 3.3550 0.5500 ;
        RECT  3.1150 -0.1800 3.2350 0.5500 ;
        RECT  2.2750 -0.1800 2.3950 0.7100 ;
        RECT  1.4350 -0.1800 1.5550 0.7100 ;
        RECT  0.5350 -0.1800 0.6550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  10.7150 1.7400 10.8350 2.7900 ;
        RECT  9.3350 1.6000 9.4550 2.7900 ;
        RECT  7.3450 1.8500 7.4650 2.7900 ;
        RECT  5.2750 2.0700 5.5150 2.1900 ;
        RECT  5.2750 2.0700 5.3950 2.7900 ;
        RECT  3.4350 2.0100 3.6750 2.1300 ;
        RECT  3.4350 2.0100 3.5550 2.7900 ;
        RECT  2.4750 2.0100 2.7150 2.1300 ;
        RECT  2.4750 2.0100 2.5950 2.7900 ;
        RECT  1.5150 2.0100 1.7550 2.1300 ;
        RECT  1.5150 2.0100 1.6350 2.7900 ;
        RECT  0.6150 2.1100 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.4600 1.5000 11.3600 1.5000 11.3600 1.8000 11.2400 1.8000 11.2400 1.6200
                 10.2150 1.6200 10.2150 1.2400 10.3350 1.2400 10.3350 1.5000 11.2400 1.5000
                 11.2400 1.3800 11.3400 1.3800 11.3400 0.5800 11.4600 0.5800 ;
        POLYGON  10.4000 0.8500 9.8550 0.8500 9.8550 1.0800 9.7400 1.0800 9.7400 1.5600 10.0950 1.5600
                 10.0950 2.2100 9.9750 2.2100 9.9750 1.6800 9.6200 1.6800 9.6200 1.4800 8.7850 1.4800
                 8.7850 1.5600 8.5850 1.5600 8.5850 2.0100 8.4650 2.0100 8.4650 1.4400 8.6650 1.4400
                 8.6650 0.8400 8.6250 0.8400 8.6250 0.6000 8.7450 0.6000 8.7450 0.7200 8.7850 0.7200
                 8.7850 1.3600 9.6200 1.3600 9.6200 0.9600 9.7350 0.9600 9.7350 0.7300 10.2800 0.7300
                 10.2800 0.5900 10.4000 0.5900 ;
        POLYGON  9.1350 0.6800 9.0150 0.6800 9.0150 0.4800 8.5050 0.4800 8.5050 0.9600 8.5450 0.9600
                 8.5450 1.3200 8.3450 1.3200 8.3450 2.1300 8.8550 2.1300 8.8550 1.6800 8.9750 1.6800
                 8.9750 2.2500 8.2250 2.2500 8.2250 1.3200 8.0050 1.3200 8.0050 1.4400 7.8850 1.4400
                 7.8850 1.2000 8.4250 1.2000 8.4250 1.0800 8.3850 1.0800 8.3850 0.3600 9.1350 0.3600 ;
        POLYGON  8.2650 1.0500 7.7650 1.0500 7.7650 1.5600 8.1050 1.5600 8.1050 2.2100 7.9850 2.2100
                 7.9850 1.6800 6.7150 1.6800 6.7150 1.8200 6.5950 1.8200 6.5950 1.4900 6.6550 1.4900
                 6.6550 0.7500 6.6350 0.7500 6.6350 0.6300 6.8750 0.6300 6.8750 0.7500 6.7750 0.7500
                 6.7750 1.5600 7.6450 1.5600 7.6450 0.9300 8.1450 0.9300 8.1450 0.6200 8.2650 0.6200 ;
        POLYGON  7.2050 0.8100 7.0850 0.8100 7.0850 0.5100 6.5150 0.5100 6.5150 1.1300 6.5350 1.1300
                 6.5350 1.3700 6.4750 1.3700 6.4750 1.9400 6.9850 1.9400 6.9850 2.0300 7.1050 2.0300
                 7.1050 2.1500 6.8650 2.1500 6.8650 2.0600 6.3550 2.0600 6.3550 1.1300 6.3950 1.1300
                 6.3950 0.5100 5.9150 0.5100 5.9150 0.9100 5.9950 0.9100 5.9950 1.1500 5.7950 1.1500
                 5.7950 0.6100 5.0350 0.6100 5.0350 0.5100 4.5550 0.5100 4.5550 0.9700 4.8150 0.9700
                 4.8150 1.0900 4.4350 1.0900 4.4350 0.3900 5.1550 0.3900 5.1550 0.4900 5.7950 0.4900
                 5.7950 0.3900 7.2050 0.3900 ;
        POLYGON  6.2750 0.7500 6.2350 0.7500 6.2350 1.9900 6.1150 1.9900 6.1150 1.3900 5.3150 1.3900
                 5.3150 1.3100 5.1750 1.3100 5.1750 1.1900 5.4350 1.1900 5.4350 1.2700 6.1150 1.2700
                 6.1150 0.7500 6.0350 0.7500 6.0350 0.6300 6.2750 0.6300 ;
        POLYGON  6.0750 2.2500 5.8350 2.2500 5.8350 1.9500 4.5550 1.9500 4.5550 2.2300 3.9050 2.2300
                 3.9050 1.8900 0.1350 1.8900 0.1350 1.7100 0.1200 1.7100 0.1200 0.7800 0.1350 0.7800
                 0.1350 0.6600 0.2550 0.6600 0.2550 0.9000 0.2400 0.9000 0.2400 1.5900 0.2550 1.5900
                 0.2550 1.7700 3.7150 1.7700 3.7150 0.9100 3.8350 0.9100 3.8350 1.7700 4.0250 1.7700
                 4.0250 2.1100 4.4350 2.1100 4.4350 1.3300 4.2150 1.3300 4.2150 1.2100 4.5550 1.2100
                 4.5550 1.8300 5.9550 1.8300 5.9550 2.1300 6.0750 2.1300 ;
        POLYGON  5.6750 1.1500 5.5550 1.1500 5.5550 1.0700 5.0550 1.0700 5.0550 1.5900 4.9750 1.5900
                 4.9750 1.7100 4.8550 1.7100 4.8550 1.4700 4.9350 1.4700 4.9350 0.8500 4.6750 0.8500
                 4.6750 0.6300 4.9150 0.6300 4.9150 0.7300 5.0550 0.7300 5.0550 0.9500 5.5550 0.9500
                 5.5550 0.9100 5.6750 0.9100 ;
        POLYGON  4.3150 1.9900 4.1950 1.9900 4.1950 1.5900 3.9750 1.5900 3.9750 0.7900 3.0950 0.7900
                 3.0950 1.1300 2.9750 1.1300 2.9750 0.6700 3.9750 0.6700 3.9750 0.5700 4.0950 0.5700
                 4.0950 1.4700 4.3150 1.4700 ;
        POLYGON  3.5150 1.3700 2.8550 1.3700 2.8550 1.5300 3.1950 1.5300 3.1950 1.6500 2.7350 1.6500
                 2.7350 1.2500 2.0750 1.2500 2.0750 1.1300 2.7350 1.1300 2.7350 0.8100 2.6950 0.8100
                 2.6950 0.5700 2.8150 0.5700 2.8150 0.6900 2.8550 0.6900 2.8550 1.2500 3.3950 1.2500
                 3.3950 0.9100 3.5150 0.9100 ;
    END
END SMDFFHQX4

MACRO SMDFFHQX2
    CLASS CORE ;
    FOREIGN SMDFFHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 0.9700 1.3800 1.6400 ;
        RECT  1.2300 0.9700 1.3800 1.4400 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8800 1.2000 7.0000 1.4400 ;
        RECT  6.4500 1.3150 7.0000 1.4350 ;
        RECT  6.4500 1.1750 6.6000 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4800 0.8850 8.6300 1.1450 ;
        RECT  8.3800 1.0250 8.5000 1.3850 ;
        END
    END SE
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.6800 1.2650 8.9200 1.3850 ;
        RECT  8.8000 0.8850 8.9200 1.3850 ;
        RECT  8.7700 0.8850 8.9200 1.1450 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1400 1.2400 10.4250 1.4700 ;
        RECT  10.1650 1.2200 10.4250 1.4700 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 0.9400 10.7150 1.0900 ;
        RECT  10.5450 0.9400 10.6650 1.1800 ;
        RECT  9.8600 0.9700 10.7150 1.0900 ;
        RECT  9.4000 1.0000 10.0450 1.1200 ;
        RECT  9.2800 1.2650 9.5200 1.3850 ;
        RECT  9.4000 1.0000 9.5200 1.3850 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6000 1.2950 0.7200 2.2100 ;
        RECT  0.3600 1.1750 0.7000 1.4350 ;
        RECT  0.5800 0.6200 0.7000 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.4200 -0.1800 10.5400 0.8200 ;
        RECT  9.1400 -0.1800 9.2600 0.6400 ;
        RECT  6.9400 -0.1800 7.0600 0.7900 ;
        RECT  4.7500 0.4900 4.9900 0.6100 ;
        RECT  4.8700 -0.1800 4.9900 0.6100 ;
        RECT  2.5300 0.5000 2.7700 0.6200 ;
        RECT  2.6500 -0.1800 2.7700 0.6200 ;
        RECT  0.9400 0.4900 1.1800 0.6100 ;
        RECT  0.9400 -0.1800 1.0600 0.6100 ;
        RECT  0.1600 -0.1800 0.2800 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.2200 1.8300 10.3400 2.7900 ;
        RECT  8.8400 1.7450 8.9600 2.7900 ;
        RECT  6.8000 1.8500 6.9200 2.7900 ;
        RECT  4.7100 2.0100 4.9500 2.1300 ;
        RECT  4.7100 2.0100 4.8300 2.7900 ;
        RECT  2.4900 1.8800 2.7300 2.0000 ;
        RECT  2.4900 1.8800 2.6100 2.7900 ;
        RECT  1.0200 1.5600 1.1400 2.7900 ;
        RECT  0.1800 1.5600 0.3000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.9600 0.8200 10.9550 0.8200 10.9550 1.7100 10.8200 1.7100 10.8200 1.8300
                 10.7000 1.8300 10.7000 1.7100 9.7200 1.7100 9.7200 1.2400 9.8400 1.2400 9.8400 1.5900
                 10.8350 1.5900 10.8350 0.7000 10.8400 0.7000 10.8400 0.5800 10.9600 0.5800 ;
        POLYGON  9.9000 0.8500 9.7400 0.8500 9.7400 0.8800 9.1600 0.8800 9.1600 1.5050 9.6000 1.5050
                 9.6000 2.2100 9.4800 2.2100 9.4800 1.6250 8.2600 1.6250 8.2600 1.6800 8.0400 1.6800
                 8.0400 2.0100 7.9200 2.0100 7.9200 1.5600 8.1400 1.5600 8.1400 0.7700 8.1200 0.7700
                 8.1200 0.6500 8.3600 0.6500 8.3600 0.7700 8.2600 0.7700 8.2600 1.5050 9.0400 1.5050
                 9.0400 0.7600 9.6200 0.7600 9.6200 0.7300 9.7800 0.7300 9.7800 0.5900 9.9000 0.5900 ;
        POLYGON  8.7400 0.7650 8.6200 0.7650 8.6200 0.5300 8.0000 0.5300 8.0000 0.8900 8.0200 0.8900
                 8.0200 1.4400 7.8000 1.4400 7.8000 2.1300 8.3600 2.1300 8.3600 1.8650 8.4800 1.8650
                 8.4800 2.2500 7.6800 2.2500 7.6800 1.4400 7.3600 1.4400 7.3600 1.2000 7.4800 1.2000
                 7.4800 1.3200 7.9000 1.3200 7.9000 1.0100 7.8800 1.0100 7.8800 0.4100 8.7400 0.4100 ;
        POLYGON  7.7600 0.7700 7.6400 0.7700 7.6400 1.0300 7.2400 1.0300 7.2400 1.5600 7.5600 1.5600
                 7.5600 2.2100 7.4400 2.2100 7.4400 1.6800 6.1900 1.6800 6.1900 1.8200 6.0700 1.8200
                 6.0700 1.4700 6.1300 1.4700 6.1300 0.7200 6.0700 0.7200 6.0700 0.6000 6.3100 0.6000
                 6.3100 0.7200 6.2500 0.7200 6.2500 1.5600 7.1200 1.5600 7.1200 0.9100 7.5200 0.9100
                 7.5200 0.6500 7.7600 0.6500 ;
        POLYGON  6.6400 0.7900 6.5200 0.7900 6.5200 0.4800 5.9500 0.4800 5.9500 1.1100 6.0100 1.1100
                 6.0100 1.3500 5.9500 1.3500 5.9500 1.9400 6.4400 1.9400 6.4400 2.0300 6.5600 2.0300
                 6.5600 2.1500 6.3200 2.1500 6.3200 2.0600 5.8300 2.0600 5.8300 0.4800 5.3500 0.4800
                 5.3500 0.8800 5.4700 0.8800 5.4700 1.1200 5.2300 1.1200 5.2300 0.8500 4.5100 0.8500
                 4.5100 0.4800 4.0300 0.4800 4.0300 0.9400 4.1500 0.9400 4.1500 1.0600 3.9100 1.0600
                 3.9100 0.3600 4.6300 0.3600 4.6300 0.7300 5.2300 0.7300 5.2300 0.3600 6.6400 0.3600 ;
        POLYGON  5.7100 1.9900 5.5900 1.9900 5.5900 1.3600 4.6300 1.3600 4.6300 1.3300 4.5100 1.3300
                 4.5100 1.2100 4.7500 1.2100 4.7500 1.2400 5.5900 1.2400 5.5900 0.7200 5.4700 0.7200
                 5.4700 0.6000 5.7100 0.6000 ;
        POLYGON  5.5100 2.2500 5.0700 2.2500 5.0700 1.8900 4.3950 1.8900 4.3950 2.2300 3.1200 2.2300
                 3.1200 1.7600 1.6200 1.7600 1.6200 1.8000 1.5000 1.8000 1.5000 1.5600 1.5400 1.5600
                 1.5400 0.6800 1.7800 0.6800 1.7800 0.8000 1.6600 0.8000 1.6600 1.6400 3.1200 1.6400
                 3.1200 1.1000 3.0300 1.1000 3.0300 0.9800 3.2700 0.9800 3.2700 1.1000 3.2400 1.1000
                 3.2400 2.1100 3.6500 2.1100 3.6500 1.1300 3.7700 1.1300 3.7700 2.1100 4.2750 2.1100
                 4.2750 1.7700 5.1900 1.7700 5.1900 2.1300 5.5100 2.1300 ;
        POLYGON  5.1100 1.0900 4.3900 1.0900 4.3900 1.6500 4.1500 1.6500 4.1500 1.5300 4.2700 1.5300
                 4.2700 0.7200 4.1500 0.7200 4.1500 0.6000 4.3900 0.6000 4.3900 0.9700 5.1100 0.9700 ;
        POLYGON  3.5300 1.9900 3.4100 1.9900 3.4100 0.7800 3.0800 0.7800 3.0800 0.8600 2.5500 0.8600
                 2.5500 1.2100 2.4300 1.2100 2.4300 0.7400 2.9600 0.7400 2.9600 0.6600 3.4100 0.6600
                 3.4100 0.5400 3.5300 0.5400 ;
        POLYGON  2.8700 1.4500 2.2900 1.4500 2.2900 1.5200 2.0100 1.5200 2.0100 1.4000 2.1700 1.4000
                 2.1700 0.5600 1.4200 0.5600 1.4200 0.8500 1.0600 0.8500 1.0600 1.1200 0.8200 1.1200
                 0.8200 0.7300 1.3000 0.7300 1.3000 0.4400 2.2900 0.4400 2.2900 1.3300 2.7500 1.3300
                 2.7500 1.1300 2.8700 1.1300 ;
    END
END SMDFFHQX2

MACRO SMDFFHQX1
    CLASS CORE ;
    FOREIGN SMDFFHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.1500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.2200 0.8950 1.4600 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.3400 0.8000 1.7250 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0950 1.2000 6.2150 1.4400 ;
        RECT  5.8700 1.2000 6.2150 1.4350 ;
        RECT  5.8700 1.1750 6.0200 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5950 0.9950 7.7600 1.4350 ;
        RECT  7.5950 0.9750 7.7150 1.4400 ;
        END
    END SE
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9000 1.0000 8.0550 1.4500 ;
        RECT  7.9350 0.9750 8.0550 1.4500 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 1.2100 9.5550 1.4650 ;
        RECT  9.2550 1.2200 9.5550 1.4500 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6750 0.9700 9.7950 1.2100 ;
        RECT  8.6450 0.9700 9.7950 1.0900 ;
        RECT  9.0050 0.9400 9.2650 1.0900 ;
        RECT  8.9150 0.9700 9.1550 1.1000 ;
        RECT  8.4150 1.0100 8.7650 1.1300 ;
        RECT  8.4150 1.0100 8.5350 1.4400 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.1500 0.1800 ;
        RECT  9.4750 -0.1800 9.5950 0.8200 ;
        RECT  8.1650 -0.1800 8.2850 0.6500 ;
        RECT  6.1750 -0.1800 6.2950 0.8000 ;
        RECT  3.9050 -0.1800 4.1450 0.3600 ;
        RECT  1.7850 0.5000 2.0250 0.6200 ;
        RECT  1.7850 -0.1800 1.9050 0.6200 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.1500 2.7900 ;
        RECT  9.3850 1.8250 9.5050 2.7900 ;
        RECT  7.9350 1.8500 8.0550 2.7900 ;
        RECT  6.0850 1.8500 6.2050 2.7900 ;
        RECT  3.9050 2.0000 4.1450 2.1200 ;
        RECT  3.9050 2.0000 4.0250 2.7900 ;
        RECT  1.9250 2.0000 2.1650 2.1200 ;
        RECT  1.9250 2.0000 2.0450 2.7900 ;
        RECT  0.5550 1.8450 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.0350 1.7050 9.9850 1.7050 9.9850 1.8250 9.8650 1.8250 9.8650 1.7050 8.8850 1.7050
                 8.8850 1.2400 9.0050 1.2400 9.0050 1.5850 9.9150 1.5850 9.9150 0.8500 9.8950 0.8500
                 9.8950 0.5800 10.0150 0.5800 10.0150 0.7300 10.0350 0.7300 ;
        POLYGON  8.9550 0.8300 8.5250 0.8300 8.5250 0.8900 8.2950 0.8900 8.2950 1.5700 8.5750 1.5700
                 8.5750 1.5600 8.6950 1.5600 8.6950 2.2100 8.5750 2.2100 8.5750 1.6900 7.3250 1.6900
                 7.3250 1.8200 7.2050 1.8200 7.2050 1.5600 7.3550 1.5600 7.3550 0.8400 7.2950 0.8400
                 7.2950 0.6000 7.4150 0.6000 7.4150 0.7200 7.4750 0.7200 7.4750 1.5700 8.1750 1.5700
                 8.1750 0.7700 8.4050 0.7700 8.4050 0.7100 8.8350 0.7100 8.8350 0.5800 8.9550 0.5800 ;
        POLYGON  7.8050 0.8400 7.6850 0.8400 7.6850 0.6000 7.5850 0.6000 7.5850 0.4800 7.1750 0.4800
                 7.1750 0.9600 7.2350 0.9600 7.2350 1.4400 7.0850 1.4400 7.0850 1.9700 7.6350 1.9700
                 7.6350 2.2100 7.5150 2.2100 7.5150 2.0900 6.9650 2.0900 6.9650 1.4400 6.5750 1.4400
                 6.5750 1.2000 6.6950 1.2000 6.6950 1.3200 7.1150 1.3200 7.1150 1.0800 7.0550 1.0800
                 7.0550 0.3600 7.7050 0.3600 7.7050 0.4800 7.8050 0.4800 ;
        POLYGON  6.9350 1.0400 6.4550 1.0400 6.4550 1.5600 6.8450 1.5600 6.8450 2.2100 6.7250 2.2100
                 6.7250 1.6800 5.4250 1.6800 5.4250 1.6400 5.3050 1.6400 5.3050 1.5200 5.4250 1.5200
                 5.4250 0.7200 5.3050 0.7200 5.3050 0.6000 5.5450 0.6000 5.5450 1.5600 6.3350 1.5600
                 6.3350 0.9200 6.8150 0.9200 6.8150 0.6200 6.9350 0.6200 ;
        POLYGON  5.8750 0.8000 5.7550 0.8000 5.7550 0.4800 5.1850 0.4800 5.1850 1.1200 5.2050 1.1200
                 5.2050 1.3600 5.1850 1.3600 5.1850 1.8000 5.7250 1.8000 5.7250 1.9100 5.8450 1.9100
                 5.8450 2.0300 5.6050 2.0300 5.6050 1.9200 5.0650 1.9200 5.0650 0.4800 4.5850 0.4800
                 4.5850 0.9200 4.7050 0.9200 4.7050 1.0400 4.4650 1.0400 4.4650 0.6000 3.6650 0.6000
                 3.6650 0.4800 3.1850 0.4800 3.1850 0.9600 3.4050 0.9600 3.4050 1.2000 3.2850 1.2000
                 3.2850 1.0800 3.0650 1.0800 3.0650 0.3600 3.7850 0.3600 3.7850 0.4800 4.4650 0.4800
                 4.4650 0.3600 5.8750 0.3600 ;
        POLYGON  4.9450 1.9800 4.8250 1.9800 4.8250 1.2800 3.7650 1.2800 3.7650 1.1600 4.8250 1.1600
                 4.8250 0.7200 4.7050 0.7200 4.7050 0.6000 4.9450 0.6000 ;
        POLYGON  4.7250 2.2400 4.3700 2.2400 4.3700 1.8800 3.1650 1.8800 3.1650 2.2200 2.3600 2.2200
                 2.3600 1.8800 1.0350 1.8800 1.0350 0.6800 1.1550 0.6800 1.1550 1.7600 2.3600 1.7600
                 2.3600 1.1000 2.2850 1.1000 2.2850 0.9800 2.5250 0.9800 2.5250 1.1000 2.4800 1.1000
                 2.4800 2.1000 3.0450 2.1000 3.0450 1.3200 2.8850 1.3200 2.8850 1.2000 3.1650 1.2000
                 3.1650 1.7600 4.4900 1.7600 4.4900 2.1200 4.7250 2.1200 ;
        POLYGON  4.3450 1.0400 3.6450 1.0400 3.6450 1.6400 3.4050 1.6400 3.4050 1.5200 3.5250 1.5200
                 3.5250 0.8400 3.3050 0.8400 3.3050 0.6000 3.5450 0.6000 3.5450 0.7200 3.6450 0.7200
                 3.6450 0.9200 4.3450 0.9200 ;
        POLYGON  2.9250 1.9800 2.8050 1.9800 2.8050 1.5600 2.6450 1.5600 2.6450 0.7800 2.2650 0.7800
                 2.2650 0.8600 1.7850 0.8600 1.7850 1.1200 1.6650 1.1200 1.6650 0.7400 2.1450 0.7400
                 2.1450 0.6600 2.6450 0.6600 2.6450 0.5400 2.7650 0.5400 2.7650 1.4400 2.9250 1.4400 ;
        POLYGON  2.1650 1.3000 2.0250 1.3000 2.0250 1.3600 1.5450 1.3600 1.5450 1.5200 1.6850 1.5200
                 1.6850 1.6400 1.4250 1.6400 1.4250 0.5600 0.9150 0.5600 0.9150 1.1000 0.5350 1.1000
                 0.5350 1.2400 0.4150 1.2400 0.4150 0.9800 0.7950 0.9800 0.7950 0.4400 1.5450 0.4400
                 1.5450 1.2400 1.9050 1.2400 1.9050 1.1800 2.1650 1.1800 ;
    END
END SMDFFHQX1

MACRO SEDFFXL
    CLASS CORE ;
    FOREIGN SEDFFXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9550 0.5000 2.0750 1.4900 ;
        RECT  1.8150 0.5000 2.0750 0.6200 ;
        RECT  1.0150 0.4200 1.9350 0.5400 ;
        RECT  1.1550 0.9800 1.2750 1.2200 ;
        RECT  0.5950 0.9800 1.2750 1.1000 ;
        RECT  0.3550 0.9700 1.1450 1.0900 ;
        RECT  0.8850 0.9400 1.1450 1.1000 ;
        RECT  1.0150 0.4200 1.1350 1.1000 ;
        RECT  0.3550 0.9700 0.4750 1.2100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2200 1.0150 1.4100 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 1.2200 4.0500 1.3400 ;
        RECT  3.9300 1.1000 4.0500 1.3400 ;
        RECT  3.5500 1.1750 3.7000 1.4350 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5800 1.0400 5.7300 1.4900 ;
        RECT  5.5900 1.0400 5.7100 1.5150 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.1450 1.0600 11.2900 1.3750 ;
        RECT  11.0900 1.1150 11.2650 1.4350 ;
        END
    END CK
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.8600 1.5900 2.9800 1.8300 ;
        RECT  2.7100 1.5900 2.9800 1.7100 ;
        RECT  2.7100 0.8850 2.8300 1.7100 ;
        RECT  2.6800 0.8850 2.8300 1.1450 ;
        RECT  2.5350 0.8850 2.8300 1.0050 ;
        RECT  2.5350 0.6000 2.6550 1.0050 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1900 1.6900 6.4500 1.8100 ;
        RECT  6.1600 1.4650 6.3100 1.7250 ;
        RECT  6.1900 0.8000 6.3100 1.8100 ;
        RECT  6.0900 0.6800 6.2100 0.9200 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  11.0100 -0.1800 11.1300 0.7000 ;
        RECT  9.0200 0.4900 9.2600 0.6100 ;
        RECT  9.1400 -0.1800 9.2600 0.6100 ;
        RECT  7.2000 0.4900 7.4400 0.6100 ;
        RECT  7.3200 -0.1800 7.4400 0.6100 ;
        RECT  5.6100 -0.1800 5.7300 0.9200 ;
        RECT  3.7300 -0.1800 3.8500 0.9200 ;
        RECT  2.0550 -0.1800 2.1750 0.3800 ;
        RECT  0.6150 -0.1800 0.7350 0.8200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  11.0100 2.0000 11.2500 2.1200 ;
        RECT  11.0100 2.0000 11.1300 2.7900 ;
        RECT  8.9000 2.2900 9.1400 2.7900 ;
        RECT  7.1800 1.6300 7.3000 2.7900 ;
        RECT  5.7300 2.1700 5.9700 2.2900 ;
        RECT  5.7300 2.1700 5.8500 2.7900 ;
        RECT  3.6700 2.2000 3.9100 2.7900 ;
        RECT  2.4950 2.2300 2.6150 2.7900 ;
        RECT  0.6150 1.7700 0.8550 1.8900 ;
        RECT  0.6150 1.7700 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.7300 1.7000 10.9700 1.7000 10.9700 1.8800 10.8000 1.8800 10.8000 2.2300
                 9.4400 2.2300 9.4400 2.1700 7.8200 2.1700 7.8200 2.0300 8.0600 2.0300 8.0600 2.0500
                 9.6800 2.0500 9.6800 2.1100 10.6800 2.1100 10.6800 1.7600 10.8500 1.7600
                 10.8500 0.8200 11.2500 0.8200 11.2500 0.7000 11.4300 0.7000 11.4300 0.4600
                 11.5500 0.4600 11.5500 0.8200 11.3700 0.8200 11.3700 0.9400 10.9700 0.9400
                 10.9700 1.5800 11.7300 1.5800 ;
        POLYGON  10.7100 1.6400 10.5600 1.6400 10.5600 1.9900 9.9600 1.9900 9.9600 1.9300 8.1800 1.9300
                 8.1800 1.3700 7.7000 1.3700 7.7000 1.2500 8.1800 1.2500 8.1800 1.2100 8.5200 1.2100
                 8.5200 1.3300 8.3000 1.3300 8.3000 1.8100 9.9600 1.8100 9.9600 1.3700 9.8400 1.3700
                 9.8400 1.2500 10.0800 1.2500 10.0800 1.8700 10.4400 1.8700 10.4400 1.5200
                 10.5900 1.5200 10.5900 0.4600 10.7100 0.4600 ;
        POLYGON  10.3200 1.7500 10.2000 1.7500 10.2000 0.4800 9.5250 0.4800 9.5250 0.8500 8.7800 0.8500
                 8.7800 0.4800 7.6800 0.4800 7.6800 0.8500 6.9600 0.8500 6.9600 0.4800 6.2850 0.4800
                 6.2850 0.5600 5.9700 0.5600 5.9700 1.7550 5.2700 1.7550 5.2700 1.8100 4.9500 1.8100
                 4.9500 0.8600 4.9100 0.8600 4.9100 0.7400 5.1500 0.7400 5.1500 0.8600 5.0700 0.8600
                 5.0700 1.6350 5.8500 1.6350 5.8500 0.4400 6.1650 0.4400 6.1650 0.3600 7.0800 0.3600
                 7.0800 0.7300 7.5600 0.7300 7.5600 0.3600 8.9000 0.3600 8.9000 0.7300 9.4050 0.7300
                 9.4050 0.3600 10.3200 0.3600 ;
        POLYGON  9.9600 1.0900 9.7200 1.0900 9.7200 1.5700 9.8400 1.5700 9.8400 1.6900 9.6000 1.6900
                 9.6000 1.4500 9.0400 1.4500 9.0400 1.3700 8.8800 1.3700 8.8800 1.2500 9.1600 1.2500
                 9.1600 1.3300 9.6000 1.3300 9.6000 0.9700 9.7200 0.9700 9.7200 0.6000 9.9600 0.6000 ;
        POLYGON  9.4000 1.2100 9.2800 1.2100 9.2800 1.1300 8.7600 1.1300 8.7600 1.6900 8.4200 1.6900
                 8.4200 1.5700 8.6400 1.5700 8.6400 1.0900 8.4200 1.0900 8.4200 0.6000 8.6600 0.6000
                 8.6600 0.9700 8.7600 0.9700 8.7600 1.0100 9.2800 1.0100 9.2800 0.9700 9.4000 0.9700 ;
        POLYGON  8.2400 0.7200 8.1200 0.7200 8.1200 1.0900 7.5800 1.0900 7.5800 1.4900 7.8800 1.4900
                 7.8800 1.5700 8.0000 1.5700 8.0000 1.6900 7.7600 1.6900 7.7600 1.6100 7.4600 1.6100
                 7.4600 1.3300 6.7400 1.3300 6.7400 1.2100 7.4600 1.2100 7.4600 0.9700 8.0000 0.9700
                 8.0000 0.6000 8.2400 0.6000 ;
        POLYGON  7.3400 1.0900 6.6200 1.0900 6.6200 1.4500 6.7800 1.4500 6.7800 1.8700 6.7700 1.8700
                 6.7700 2.0500 6.3300 2.0500 6.3300 2.2500 6.0900 2.2500 6.0900 2.0500 5.4450 2.0500
                 5.4450 2.1100 4.2650 2.1100 4.2650 2.0800 3.3500 2.0800 3.3500 1.9600 4.3850 1.9600
                 4.3850 1.9900 5.3250 1.9900 5.3250 1.9300 6.6500 1.9300 6.6500 1.7500 6.6600 1.7500
                 6.6600 1.5700 6.5000 1.5700 6.5000 0.6000 6.8400 0.6000 6.8400 0.7200 6.6200 0.7200
                 6.6200 0.9700 7.3400 0.9700 ;
        POLYGON  5.4300 1.4700 5.1900 1.4700 5.1900 1.3500 5.2700 1.3500 5.2700 0.6200 4.2700 0.6200
                 4.2700 0.8000 4.2900 0.8000 4.2900 1.4800 4.3900 1.4800 4.3900 1.6000 4.1500 1.6000
                 4.1500 1.4800 4.1700 1.4800 4.1700 0.9200 4.1500 0.9200 4.1500 0.5000 4.7500 0.5000
                 4.7500 0.4000 4.9900 0.4000 4.9900 0.5000 5.3900 0.5000 5.3900 1.3500 5.4300 1.3500 ;
        POLYGON  4.7900 1.8700 4.6700 1.8700 4.6700 1.8400 3.2200 1.8400 3.2200 2.0700 1.7350 2.0700
                 1.7350 1.8300 1.7150 1.8300 1.7150 0.8600 1.2550 0.8600 1.2550 0.6600 1.4950 0.6600
                 1.4950 0.7400 1.8350 0.7400 1.8350 1.7100 1.8550 1.7100 1.8550 1.9500 3.1000 1.9500
                 3.1000 1.7200 4.6700 1.7200 4.6700 0.8600 4.4900 0.8600 4.4900 0.7400 4.7900 0.7400 ;
        POLYGON  3.4300 1.6000 3.1900 1.6000 3.1900 1.4800 3.3100 1.4800 3.3100 0.6800 2.8250 0.6800
                 2.8250 0.4800 2.4150 0.4800 2.4150 1.1600 2.2950 1.1600 2.2950 0.3600 2.9450 0.3600
                 2.9450 0.5600 3.4300 0.5600 ;
        POLYGON  1.5950 1.6500 0.3750 1.6500 0.3750 1.8300 0.2550 1.8300 0.2550 1.7100 0.1150 1.7100
                 0.1150 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000 0.2550 0.8400 0.2350 0.8400
                 0.2350 1.5300 1.4750 1.5300 1.4750 1.2500 1.5950 1.2500 ;
    END
END SEDFFXL

MACRO SEDFFX4
    CLASS CORE ;
    FOREIGN SEDFFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.5000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4050 1.5000 1.5250 2.1500 ;
        RECT  1.4050 0.6800 1.5250 1.0250 ;
        RECT  1.3850 0.9050 1.5050 1.6200 ;
        RECT  0.5650 1.0250 1.5050 1.1450 ;
        RECT  0.5650 0.8850 0.8000 1.1450 ;
        RECT  0.5650 0.6800 0.6850 2.1500 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8450 1.2300 8.1050 1.5000 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1350 0.8950 8.3950 1.1100 ;
        RECT  8.2450 0.8950 8.3650 1.2750 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1850 1.0900 10.3700 1.5050 ;
        RECT  10.1850 1.0900 10.3050 1.5200 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.3700 1.4300 13.5850 1.6700 ;
        RECT  13.3250 1.4650 13.5600 1.7250 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.1300 1.1250 13.9850 1.2450 ;
        RECT  13.7000 0.8850 13.8500 1.2450 ;
        RECT  12.6650 1.2250 13.2500 1.3450 ;
        RECT  12.6650 1.2250 12.7850 1.7500 ;
        END
    END E
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0900 0.8500 11.9050 0.9700 ;
        RECT  11.7850 0.6800 11.9050 0.9700 ;
        RECT  11.5850 1.6200 11.8250 1.7400 ;
        RECT  11.0900 1.5000 11.7050 1.6200 ;
        RECT  11.0900 1.4650 11.2400 1.7250 ;
        RECT  10.6250 1.6200 11.2100 1.7400 ;
        RECT  11.0900 0.8000 11.2100 1.7400 ;
        RECT  10.9450 0.8000 11.2100 0.9200 ;
        RECT  10.9450 0.6800 11.0650 0.9200 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.5000 0.1800 ;
        RECT  13.5850 -0.1800 13.7050 0.7650 ;
        RECT  12.2050 -0.1800 12.3250 0.7300 ;
        RECT  11.3650 -0.1800 11.4850 0.7300 ;
        RECT  10.5250 -0.1800 10.6450 0.7300 ;
        RECT  8.2250 0.4150 8.4650 0.5350 ;
        RECT  8.3450 -0.1800 8.4650 0.5350 ;
        RECT  6.7900 -0.1800 6.9100 0.7300 ;
        RECT  4.4450 0.6100 4.6850 0.7300 ;
        RECT  4.5650 -0.1800 4.6850 0.7300 ;
        RECT  2.7250 -0.1800 2.8450 0.8200 ;
        RECT  1.8250 -0.1800 1.9450 0.7300 ;
        RECT  0.9850 -0.1800 1.1050 0.7300 ;
        RECT  0.1450 -0.1800 0.2650 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.5000 2.7900 ;
        RECT  13.6250 2.0850 13.7450 2.7900 ;
        RECT  12.0650 2.1000 12.3050 2.2200 ;
        RECT  12.0650 2.1000 12.1850 2.7900 ;
        RECT  11.1050 2.1000 11.3450 2.2200 ;
        RECT  11.1050 2.1000 11.2250 2.7900 ;
        RECT  10.1450 2.1000 10.3850 2.2200 ;
        RECT  10.1450 2.1000 10.2650 2.7900 ;
        RECT  8.2350 1.8600 8.3550 2.7900 ;
        RECT  6.6450 1.8800 6.7650 2.7900 ;
        RECT  6.5250 1.8800 6.7650 2.0000 ;
        RECT  4.6250 1.8100 4.7450 2.7900 ;
        RECT  4.5050 1.8100 4.7450 1.9300 ;
        RECT  2.7250 2.0200 2.8450 2.7900 ;
        RECT  1.8250 1.6300 1.9450 2.7900 ;
        RECT  0.9850 1.5000 1.1050 2.7900 ;
        RECT  0.1450 1.5000 0.2650 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.2250 2.0900 14.1050 2.0900 14.1050 1.9650 13.0650 1.9650 13.0650 1.5300
                 13.1850 1.5300 13.1850 1.8450 14.1050 1.8450 14.1050 1.0050 14.0050 1.0050
                 14.0050 0.5250 14.1250 0.5250 14.1250 0.8850 14.2250 0.8850 ;
        POLYGON  13.0650 0.9700 12.5450 0.9700 12.5450 1.8700 12.9450 1.8700 12.9450 2.1100
                 12.8250 2.1100 12.8250 1.9900 12.4250 1.9900 12.4250 1.9800 9.2950 1.9800
                 9.2950 1.3800 9.5850 1.3800 9.5850 0.8600 9.5050 0.8600 9.5050 0.6000 9.6250 0.6000
                 9.6250 0.7400 9.7050 0.7400 9.7050 1.5000 9.4150 1.5000 9.4150 1.8600 12.4250 1.8600
                 12.4250 0.8500 12.9450 0.8500 12.9450 0.5250 13.0650 0.5250 ;
        POLYGON  10.7850 1.2400 10.6650 1.2400 10.6650 1.0900 10.5500 1.0900 10.5500 0.9700
                 10.2850 0.9700 10.2850 0.5600 9.8400 0.5600 9.8400 0.4800 8.9000 0.4800 8.9000 0.7750
                 7.9850 0.7750 7.9850 0.4800 7.3300 0.4800 7.3300 0.8000 7.4850 0.8000 7.4850 1.7700
                 7.3650 1.7700 7.3650 0.9200 7.2100 0.9200 7.2100 0.3600 8.1050 0.3600 8.1050 0.6550
                 8.7800 0.6550 8.7800 0.3600 9.9600 0.3600 9.9600 0.4400 10.4050 0.4400 10.4050 0.8500
                 10.6700 0.8500 10.6700 0.9700 10.7850 0.9700 ;
        POLYGON  10.1650 0.9200 9.9450 0.9200 9.9450 1.7400 9.6650 1.7400 9.6650 1.6200 9.8250 1.6200
                 9.8250 0.8000 10.0450 0.8000 10.0450 0.6800 10.1650 0.6800 ;
        POLYGON  9.4650 1.2600 8.9650 1.2600 8.9650 1.6000 8.7250 1.6000 8.7250 1.4800 8.8450 1.4800
                 8.8450 1.1400 9.3450 1.1400 9.3450 0.9800 9.4650 0.9800 ;
        POLYGON  9.2050 1.0200 8.6350 1.0200 8.6350 1.3600 8.6050 1.3600 8.6050 1.8000 9.0550 1.8000
                 9.0550 1.9200 8.4850 1.9200 8.4850 1.7400 8.1150 1.7400 8.1150 2.2500 6.8850 2.2500
                 6.8850 1.7600 5.7450 1.7600 5.7450 1.8700 5.6250 1.8700 5.6250 1.6100 5.8050 1.6100
                 5.8050 0.8600 5.7450 0.8600 5.7450 0.6200 5.8650 0.6200 5.8650 0.7400 5.9250 0.7400
                 5.9250 1.6400 7.0050 1.6400 7.0050 2.1300 7.9950 2.1300 7.9950 1.6200 8.4850 1.6200
                 8.4850 1.2400 8.5150 1.2400 8.5150 0.9000 9.0850 0.9000 9.0850 0.6000 9.2050 0.6000 ;
        POLYGON  7.8750 2.0100 7.1250 2.0100 7.1250 1.2000 6.3250 1.2000 6.3250 1.0800 7.2450 1.0800
                 7.2450 1.8900 7.6050 1.8900 7.6050 0.9900 7.7450 0.9900 7.7450 0.6000 7.8650 0.6000
                 7.8650 1.1100 7.7250 1.1100 7.7250 1.7400 7.8750 1.7400 ;
        POLYGON  6.4300 0.9200 6.2050 0.9200 6.2050 1.4000 6.2850 1.4000 6.2850 1.5200 6.0450 1.5200
                 6.0450 1.4000 6.0850 1.4000 6.0850 0.8000 6.3100 0.8000 6.3100 0.6800 6.0450 0.6800
                 6.0450 0.5000 5.6250 0.5000 5.6250 1.3700 5.6850 1.3700 5.6850 1.4900 5.4450 1.4900
                 5.4450 1.3700 5.5050 1.3700 5.5050 0.5000 4.9250 0.5000 4.9250 0.9700 4.2050 0.9700
                 4.2050 0.5000 3.3650 0.5000 3.3650 1.1800 3.3850 1.1800 3.3850 1.4200 3.2450 1.4200
                 3.2450 0.3800 3.7650 0.3800 3.7650 0.3600 4.0050 0.3600 4.0050 0.3800 4.3250 0.3800
                 4.3250 0.8500 4.8050 0.8500 4.8050 0.3800 5.0050 0.3800 5.0050 0.3600 5.2450 0.3600
                 5.2450 0.3800 6.1650 0.3800 6.1650 0.5600 6.4300 0.5600 ;
        POLYGON  6.4050 2.2000 5.3950 2.2000 5.3950 2.1100 4.8650 2.1100 4.8650 1.6900 4.3850 1.6900
                 4.3850 2.1100 3.7450 2.1100 3.7450 2.0500 3.2450 2.0500 3.2450 2.2500 3.0050 2.2500
                 3.0050 1.9000 2.3650 1.9000 2.3650 2.1500 2.2450 2.1500 2.2450 1.7500 2.2050 1.7500
                 2.2050 1.3600 1.6250 1.3600 1.6250 1.2400 2.2050 1.2400 2.2050 0.8000 2.3050 0.8000
                 2.3050 0.6800 2.4250 0.6800 2.4250 0.9200 2.3250 0.9200 2.3250 1.6300 2.3650 1.6300
                 2.3650 1.7800 3.1250 1.7800 3.1250 1.9300 3.8650 1.9300 3.8650 1.9900 4.2650 1.9900
                 4.2650 1.5700 4.9850 1.5700 4.9850 1.9900 5.5150 1.9900 5.5150 2.0800 6.4050 2.0800 ;
        POLYGON  5.3850 0.8000 5.2650 0.8000 5.2650 1.6300 5.3250 1.6300 5.3250 1.8700 5.2050 1.8700
                 5.2050 1.7500 5.1450 1.7500 5.1450 1.2100 4.2250 1.2100 4.2250 1.0900 5.1450 1.0900
                 5.1450 0.6800 5.3850 0.6800 ;
        POLYGON  4.9050 1.4500 4.1050 1.4500 4.1050 1.8700 3.9850 1.8700 3.9850 1.2100 3.9650 1.2100
                 3.9650 0.6200 4.0850 0.6200 4.0850 1.0900 4.1050 1.0900 4.1050 1.3300 4.9050 1.3300 ;
        POLYGON  3.7450 1.8100 3.5050 1.8100 3.5050 1.6600 3.0050 1.6600 3.0050 1.4700 2.4450 1.4700
                 2.4450 1.3500 3.1250 1.3500 3.1250 1.5400 3.5050 1.5400 3.5050 0.8000 3.4850 0.8000
                 3.4850 0.6800 3.7250 0.6800 3.7250 0.8000 3.6250 0.8000 3.6250 1.6900 3.7450 1.6900 ;
    END
END SEDFFX4

MACRO SEDFFX2
    CLASS CORE ;
    FOREIGN SEDFFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.7600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9050 1.2800 7.0250 1.5200 ;
        RECT  6.7400 1.2800 7.0250 1.4350 ;
        RECT  6.7400 1.1750 6.8900 1.4350 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.2300 7.5250 1.4450 ;
        RECT  7.3250 1.2300 7.4450 1.6400 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 1.1800 9.5550 1.4500 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6150 1.2100 11.9150 1.4250 ;
        RECT  11.6150 1.2100 11.8750 1.4500 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 1.2300 12.4550 1.3800 ;
        RECT  12.1650 1.2100 12.3150 1.3300 ;
        RECT  12.1650 0.9700 12.2850 1.3300 ;
        RECT  11.0450 0.9700 12.2850 1.0900 ;
        RECT  11.0450 0.9700 11.4950 1.1700 ;
        RECT  11.0450 0.9700 11.1650 1.7700 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6800 0.6750 1.9900 ;
        RECT  0.3600 0.8850 0.6750 1.1450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.9450 1.4650 10.1850 1.7400 ;
        RECT  10.0650 0.6700 10.1850 1.7400 ;
        RECT  9.9300 1.4650 10.1850 1.7250 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.7600 0.1800 ;
        RECT  11.8150 0.7300 12.0550 0.8500 ;
        RECT  11.8150 -0.1800 11.9350 0.8500 ;
        RECT  10.5450 -0.1800 10.6650 0.3900 ;
        RECT  9.5850 0.5400 9.8250 0.6600 ;
        RECT  9.7050 -0.1800 9.8250 0.6600 ;
        RECT  7.1650 -0.1800 7.2850 0.8000 ;
        RECT  5.5400 -0.1800 5.6600 0.9000 ;
        RECT  3.4000 0.6100 3.6400 0.7300 ;
        RECT  3.5200 -0.1800 3.6400 0.7300 ;
        RECT  1.8000 -0.1800 1.9200 0.5300 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.7600 2.7900 ;
        RECT  11.9050 1.9700 12.0250 2.7900 ;
        RECT  10.4250 2.1000 10.6650 2.2200 ;
        RECT  10.4250 2.1000 10.5450 2.7900 ;
        RECT  9.4650 2.1000 9.7050 2.2200 ;
        RECT  9.4650 2.1000 9.5850 2.7900 ;
        RECT  7.2650 2.2400 7.5050 2.7900 ;
        RECT  5.5400 1.8800 5.6600 2.7900 ;
        RECT  5.4200 1.8800 5.6600 2.0000 ;
        RECT  3.5200 1.8100 3.6400 2.7900 ;
        RECT  3.4000 1.8100 3.6400 1.9300 ;
        RECT  1.6400 2.0100 1.7600 2.7900 ;
        RECT  1.0350 2.1400 1.1550 2.7900 ;
        RECT  0.1350 1.3400 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.6950 1.9700 12.4450 1.9700 12.4450 2.0900 12.3250 2.0900 12.3250 1.8500
                 12.5750 1.8500 12.5750 1.6900 11.3450 1.6900 11.3450 1.5700 12.5750 1.5700
                 12.5750 0.8500 12.2350 0.8500 12.2350 0.7300 12.6950 0.7300 ;
        POLYGON  11.4150 0.8500 10.9250 0.8500 10.9250 1.9100 11.3650 1.9100 11.3650 2.0300
                 10.8050 2.0300 10.8050 1.9800 8.4450 1.9800 8.4450 1.6200 8.7450 1.6200 8.7450 0.7400
                 8.1650 0.7400 8.1650 0.6200 8.8650 0.6200 8.8650 1.7400 8.5650 1.7400 8.5650 1.8600
                 10.8050 1.8600 10.8050 0.7300 11.4150 0.7300 ;
        POLYGON  9.9050 1.2300 9.7850 1.2300 9.7850 0.9000 9.3450 0.9000 9.3450 0.5000 7.5250 0.5000
                 7.5250 1.0400 6.9250 1.0400 6.9250 0.5000 6.2500 0.5000 6.2500 0.6600 6.0800 0.6600
                 6.0800 0.9000 6.3800 0.9000 6.3800 1.5800 6.2600 1.5800 6.2600 1.0200 5.9600 1.0200
                 5.9600 0.5400 6.1300 0.5400 6.1300 0.3800 7.0450 0.3800 7.0450 0.9200 7.4050 0.9200
                 7.4050 0.3800 9.4650 0.3800 9.4650 0.7800 9.9050 0.7800 ;
        POLYGON  9.2250 0.7400 9.1050 0.7400 9.1050 0.9400 9.2250 0.9400 9.2250 1.0600 9.1050 1.0600
                 9.1050 1.6200 9.2250 1.6200 9.2250 1.7400 8.9850 1.7400 8.9850 0.6200 9.2250 0.6200 ;
        POLYGON  8.6250 1.5000 7.8850 1.5000 7.8850 1.3800 8.5050 1.3800 8.5050 0.9000 8.6250 0.9000 ;
        POLYGON  8.1450 1.8800 8.0250 1.8800 8.0250 1.7600 7.7650 1.7600 7.7650 1.8800 7.2350 1.8800
                 7.2350 2.1200 6.3200 2.1200 6.3200 2.0600 5.7800 2.0600 5.7800 1.7600 4.8400 1.7600
                 4.8400 1.7700 4.7000 1.7700 4.7000 1.8900 4.5800 1.8900 4.5800 1.6500 4.7000 1.6500
                 4.7000 0.6200 4.8200 0.6200 4.8200 1.6400 5.9000 1.6400 5.9000 1.9400 6.4400 1.9400
                 6.4400 2.0000 7.1150 2.0000 7.1150 1.7600 7.6450 1.7600 7.6450 1.1400 7.7450 1.1400
                 7.7450 0.6200 7.9850 0.6200 7.9850 0.7400 7.8650 0.7400 7.8650 1.2600 7.7650 1.2600
                 7.7650 1.6400 8.1450 1.6400 ;
        POLYGON  6.9650 1.8800 6.8450 1.8800 6.8450 1.8200 6.0200 1.8200 6.0200 1.5200 5.8100 1.5200
                 5.8100 1.2600 5.2800 1.2600 5.2800 1.0200 5.4000 1.0200 5.4000 1.1400 5.9300 1.1400
                 5.9300 1.4000 6.1400 1.4000 6.1400 1.7000 6.5000 1.7000 6.5000 0.6200 6.8050 0.6200
                 6.8050 0.7400 6.6200 0.7400 6.6200 1.6400 6.9650 1.6400 ;
        POLYGON  5.3000 2.2000 3.7600 2.2000 3.7600 1.6900 3.2800 1.6900 3.2800 2.1100 2.1600 2.1100
                 2.1600 2.2500 1.9200 2.2500 1.9200 2.1300 2.0400 2.1300 2.0400 1.8900 1.6600 1.8900
                 1.6600 1.8400 1.3950 1.8400 1.3950 1.4600 1.2150 1.4600 1.2150 1.2000 0.7950 1.2000
                 0.7950 1.0800 1.2150 1.0800 1.2150 0.7400 1.6350 0.7400 1.6350 0.8600 1.3350 0.8600
                 1.3350 1.3400 1.5150 1.3400 1.5150 1.7200 1.7800 1.7200 1.7800 1.7700 2.1600 1.7700
                 2.1600 1.9900 3.1600 1.9900 3.1600 1.5700 3.8800 1.5700 3.8800 2.0800 5.3000 2.0800 ;
        POLYGON  5.2400 0.9000 5.1600 0.9000 5.1600 1.4000 5.1800 1.4000 5.1800 1.5200 4.9400 1.5200
                 4.9400 1.4000 5.0400 1.4000 5.0400 0.7800 5.1200 0.7800 5.1200 0.6600 4.9400 0.6600
                 4.9400 0.5000 4.5800 0.5000 4.5800 1.0400 4.5600 1.0400 4.5600 1.5300 4.4400 1.5300
                 4.4400 0.9200 4.4600 0.9200 4.4600 0.5000 3.8800 0.5000 3.8800 0.9700 3.1600 0.9700
                 3.1600 0.5000 2.3200 0.5000 2.3200 1.2900 2.4000 1.2900 2.4000 1.4100 2.1600 1.4100
                 2.1600 1.2900 2.2000 1.2900 2.2000 0.3800 2.6100 0.3800 2.6100 0.3600 2.8500 0.3600
                 2.8500 0.3800 3.2800 0.3800 3.2800 0.8500 3.7600 0.8500 3.7600 0.3800 3.9600 0.3800
                 3.9600 0.3600 4.2000 0.3600 4.2000 0.3800 5.0600 0.3800 5.0600 0.5400 5.2400 0.5400 ;
        POLYGON  4.3400 0.8000 4.2200 0.8000 4.2200 1.6300 4.2800 1.6300 4.2800 1.8700 4.1600 1.8700
                 4.1600 1.7500 4.1000 1.7500 4.1000 1.2100 3.1800 1.2100 3.1800 1.0900 4.1000 1.0900
                 4.1000 0.6800 4.3400 0.6800 ;
        POLYGON  3.8400 1.4500 3.0400 1.4500 3.0400 1.8700 2.9200 1.8700 2.9200 0.6200 3.0400 0.6200
                 3.0400 1.3300 3.8400 1.3300 ;
        POLYGON  2.6800 0.8000 2.6400 0.8000 2.6400 1.6900 2.6800 1.6900 2.6800 1.8100 2.4400 1.8100
                 2.4400 1.6500 1.9000 1.6500 1.9000 1.2000 1.4550 1.2000 1.4550 1.0800 2.0200 1.0800
                 2.0200 1.5300 2.5200 1.5300 2.5200 0.8000 2.4400 0.8000 2.4400 0.6800 2.6800 0.6800 ;
    END
END SEDFFX2

MACRO SEDFFX1
    CLASS CORE ;
    FOREIGN SEDFFX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0850 0.5000 2.2050 1.4900 ;
        RECT  1.9450 0.5000 2.2050 0.6200 ;
        RECT  1.1650 0.4200 2.0650 0.5400 ;
        RECT  1.2650 0.9800 1.3850 1.2200 ;
        RECT  1.1650 0.4200 1.2850 1.1000 ;
        RECT  0.5350 0.9800 1.3850 1.1000 ;
        RECT  0.3050 1.2300 0.6550 1.3800 ;
        RECT  0.5350 0.9400 0.6550 1.3800 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.2200 1.1450 1.4100 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9400 1.0550 4.0850 1.2950 ;
        RECT  3.8400 1.1750 4.0100 1.4350 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5800 0.8100 5.7300 1.2650 ;
        RECT  5.5900 0.8100 5.7100 1.5300 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0900 1.0850 11.3100 1.4350 ;
        END
    END CK
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7100 1.5700 3.2300 1.6900 ;
        RECT  2.7100 0.7200 2.8300 1.6900 ;
        RECT  2.6650 0.6000 2.7850 0.8400 ;
        RECT  2.6800 1.1750 2.8300 1.4350 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3300 1.6200 6.5700 1.8650 ;
        RECT  6.3300 0.7600 6.4500 1.8650 ;
        RECT  6.1050 0.7600 6.4500 1.0900 ;
        RECT  6.1050 0.6400 6.2250 1.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  11.0300 -0.1800 11.1500 0.7250 ;
        RECT  9.0400 0.3100 9.2800 0.4300 ;
        RECT  9.0400 -0.1800 9.1600 0.4300 ;
        RECT  7.3000 0.4500 7.5400 0.5700 ;
        RECT  7.3000 -0.1800 7.4200 0.5700 ;
        RECT  5.6250 -0.1800 5.7450 0.6900 ;
        RECT  3.6950 -0.1800 3.8150 0.9200 ;
        RECT  2.1850 -0.1800 2.3050 0.3800 ;
        RECT  0.7250 0.6600 0.9650 0.7800 ;
        RECT  0.8450 -0.1800 0.9650 0.7800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  11.0900 1.7950 11.2100 2.7900 ;
        RECT  8.9200 2.2900 9.1600 2.7900 ;
        RECT  7.2600 2.1500 7.3800 2.7900 ;
        RECT  5.8500 2.2250 6.0900 2.7900 ;
        RECT  3.8600 2.2900 4.1000 2.7900 ;
        RECT  2.5700 2.2300 2.6900 2.7900 ;
        RECT  0.7250 1.7700 0.9650 1.8900 ;
        RECT  0.7250 1.7700 0.8450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6900 1.8550 11.4500 1.8550 11.4500 1.6750 10.9700 1.6750 10.9700 2.2300
                 9.4600 2.2300 9.4600 2.1700 8.1600 2.1700 8.1600 2.0500 9.7000 2.0500 9.7000 2.1100
                 10.8500 2.1100 10.8500 0.8450 11.2700 0.8450 11.2700 0.6050 11.4500 0.6050
                 11.4500 0.4850 11.5700 0.4850 11.5700 0.7250 11.3900 0.7250 11.3900 0.9650
                 10.9700 0.9650 10.9700 1.5550 11.5700 1.5550 11.5700 1.7350 11.6900 1.7350 ;
        POLYGON  10.7300 1.9900 9.9800 1.9900 9.9800 1.9300 8.2600 1.9300 8.2600 1.2900 7.9200 1.2900
                 7.9200 1.4100 7.8000 1.4100 7.8000 1.1700 8.2600 1.1700 8.2600 1.0300 8.5400 1.0300
                 8.5400 1.1500 8.3800 1.1500 8.3800 1.8100 9.9800 1.8100 9.9800 1.4100 9.9400 1.4100
                 9.9400 1.1700 10.0600 1.1700 10.0600 1.2900 10.1000 1.2900 10.1000 1.8700
                 10.6100 1.8700 10.6100 0.4850 10.7300 0.4850 ;
        POLYGON  10.3400 1.7500 10.2200 1.7500 10.2200 0.4800 9.5450 0.4800 9.5450 0.6700 8.8000 0.6700
                 8.8000 0.4800 7.7800 0.4800 7.7800 0.8100 7.0600 0.8100 7.0600 0.4800 5.9850 0.4800
                 5.9850 1.1000 5.9700 1.1000 5.9700 1.8650 5.3300 1.8650 5.3300 1.9850 5.2100 1.9850
                 5.2100 1.8650 5.1000 1.8650 5.1000 0.8800 4.9250 0.8800 4.9250 0.6400 5.0450 0.6400
                 5.0450 0.7600 5.2200 0.7600 5.2200 1.7450 5.8500 1.7450 5.8500 0.9800 5.8650 0.9800
                 5.8650 0.3600 7.1800 0.3600 7.1800 0.6900 7.6600 0.6900 7.6600 0.3600 8.9200 0.3600
                 8.9200 0.5500 9.4250 0.5500 9.4250 0.3600 10.3400 0.3600 ;
        POLYGON  9.9800 0.7200 9.8200 0.7200 9.8200 1.5700 9.8600 1.5700 9.8600 1.6900 9.6200 1.6900
                 9.6200 1.5700 9.7000 1.5700 9.7000 1.3700 8.9000 1.3700 8.9000 1.2500 9.7000 1.2500
                 9.7000 0.6000 9.9800 0.6000 ;
        POLYGON  9.4200 1.1300 9.3000 1.1300 9.3000 1.0300 8.7800 1.0300 8.7800 1.6900 8.5000 1.6900
                 8.5000 1.5700 8.6600 1.5700 8.6600 0.9100 8.4400 0.9100 8.4400 0.6000 8.6800 0.6000
                 8.6800 0.7900 8.7800 0.7900 8.7800 0.9100 9.3000 0.9100 9.3000 0.8900 9.4200 0.8900 ;
        POLYGON  8.2600 0.7200 8.0200 0.7200 8.0200 1.0500 7.6800 1.0500 7.6800 1.5300 8.0200 1.5300
                 8.0200 1.5700 8.1400 1.5700 8.1400 1.6900 7.9000 1.6900 7.9000 1.6500 7.5600 1.6500
                 7.5600 1.3700 6.9800 1.3700 6.9800 1.2500 7.5600 1.2500 7.5600 0.9300 7.9000 0.9300
                 7.9000 0.6000 8.2600 0.6000 ;
        POLYGON  7.4400 1.0500 6.8600 1.0500 6.8600 1.6300 6.9000 1.6300 6.9000 2.1050 5.7300 2.1050
                 5.7300 2.2250 4.4550 2.2250 4.4550 2.1700 3.5400 2.1700 3.5400 2.0500 4.5750 2.0500
                 4.5750 2.1050 5.6100 2.1050 5.6100 1.9850 6.0900 1.9850 6.0900 1.2200 6.2100 1.2200
                 6.2100 1.9850 6.7800 1.9850 6.7800 1.7500 6.7400 1.7500 6.7400 0.7200 6.7000 0.7200
                 6.7000 0.6000 6.9400 0.6000 6.9400 0.7200 6.8600 0.7200 6.8600 0.9300 7.4400 0.9300 ;
        POLYGON  5.4700 1.6250 5.3500 1.6250 5.3500 1.5050 5.3400 1.5050 5.3400 0.5200 4.2350 0.5200
                 4.2350 0.8000 4.3250 0.8000 4.3250 1.4500 4.5200 1.4500 4.5200 1.6900 4.4000 1.6900
                 4.4000 1.5700 4.2050 1.5700 4.2050 0.9200 4.1150 0.9200 4.1150 0.4000 4.7050 0.4000
                 4.7050 0.3600 4.9450 0.3600 4.9450 0.4000 5.4600 0.4000 5.4600 1.3850 5.4700 1.3850 ;
        POLYGON  4.9100 1.9450 4.7900 1.9450 4.7900 1.9300 1.8850 1.9300 1.8850 1.7300 1.8450 1.7300
                 1.8450 0.8600 1.4050 0.8600 1.4050 0.6600 1.6450 0.6600 1.6450 0.7400 1.9650 0.7400
                 1.9650 1.6100 2.0050 1.6100 2.0050 1.8100 4.6850 1.8100 4.6850 0.8200 4.4450 0.8200
                 4.4450 0.7000 4.8050 0.7000 4.8050 1.7050 4.9100 1.7050 ;
        POLYGON  3.5600 1.6900 3.4400 1.6900 3.4400 0.9200 3.2750 0.9200 3.2750 0.6800 3.0100 0.6800
                 3.0100 0.4800 2.5450 0.4800 2.5450 1.1600 2.4250 1.1600 2.4250 0.3600 3.1300 0.3600
                 3.1300 0.5600 3.3950 0.5600 3.3950 0.8000 3.5600 0.8000 ;
        POLYGON  1.7250 1.6500 0.4850 1.6500 0.4850 1.8300 0.3650 1.8300 0.3650 1.7100 0.0650 1.7100
                 0.0650 0.9900 0.2950 0.9900 0.2950 0.6000 0.4150 0.6000 0.4150 1.1100 0.1850 1.1100
                 0.1850 1.5300 1.6050 1.5300 1.6050 1.2700 1.7250 1.2700 ;
    END
END SEDFFX1

MACRO SEDFFTRXL
    CLASS CORE ;
    FOREIGN SEDFFTRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.2100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8150 1.1500 6.0750 1.3800 ;
        RECT  5.8650 1.0400 5.9850 1.4500 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0450 0.9400 8.1650 1.2000 ;
        RECT  6.9050 0.9400 8.1650 1.0600 ;
        RECT  6.9050 0.9400 7.0250 1.3300 ;
        RECT  6.6850 1.2300 6.9450 1.3800 ;
        RECT  6.8250 1.2100 7.0250 1.3300 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.1800 7.5250 1.4500 ;
        END
    END SI
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.8650 1.3700 10.1050 1.5350 ;
        RECT  9.9300 1.3700 10.0800 1.7400 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.0850 1.1800 13.0500 1.3000 ;
        RECT  12.4850 1.1800 12.7450 1.3800 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.4100 1.1700 13.6950 1.2900 ;
        RECT  13.5750 1.0450 13.6950 1.2900 ;
        RECT  13.4100 1.1700 13.5600 1.4350 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 0.6800 0.2650 0.9400 ;
        RECT  0.1350 0.8200 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3850 0.6200 9.5050 1.4350 ;
        RECT  9.2050 1.5100 9.4750 1.6300 ;
        RECT  9.3500 1.1750 9.4750 1.6300 ;
        RECT  9.2050 1.5100 9.3250 1.7500 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.2100 0.1800 ;
        RECT  13.4350 -0.1800 13.5550 0.9200 ;
        RECT  11.9250 0.4600 12.1650 0.5800 ;
        RECT  11.9250 -0.1800 12.0450 0.5800 ;
        RECT  11.4350 0.4300 11.6750 0.5500 ;
        RECT  11.4350 -0.1800 11.5550 0.5500 ;
        RECT  10.3150 0.6000 10.5550 0.7200 ;
        RECT  10.4350 -0.1800 10.5550 0.7200 ;
        RECT  8.9050 -0.1800 9.0250 0.8150 ;
        RECT  7.0850 0.4600 7.3250 0.5800 ;
        RECT  7.0850 -0.1800 7.2050 0.5800 ;
        RECT  5.7250 -0.1800 5.8450 0.6800 ;
        RECT  3.6150 0.6100 3.8550 0.7300 ;
        RECT  3.7350 -0.1800 3.8550 0.7300 ;
        RECT  1.9150 -0.1800 2.0350 0.8600 ;
        RECT  0.5650 -0.1800 0.6850 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.2100 2.7900 ;
        RECT  13.4950 2.0800 13.6150 2.7900 ;
        RECT  10.0750 2.2300 10.1950 2.7900 ;
        RECT  8.6650 2.2500 8.9050 2.7900 ;
        RECT  7.0850 2.2900 7.3250 2.7900 ;
        RECT  5.6350 2.2900 5.8750 2.7900 ;
        RECT  3.7350 1.8100 3.8550 2.7900 ;
        RECT  3.6150 1.8100 3.8550 1.9300 ;
        RECT  1.8550 1.9400 1.9750 2.7900 ;
        RECT  0.5550 2.1600 0.7950 2.2800 ;
        RECT  0.5550 2.1600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.0750 1.9200 13.2800 1.9200 13.2800 2.1800 12.4250 2.1800 12.4250 2.0600
                 13.1600 2.0600 13.1600 1.8000 13.9550 1.8000 13.9550 1.6800 13.8550 1.6800
                 13.8550 0.6800 13.9750 0.6800 13.9750 1.5600 14.0750 1.5600 ;
        POLYGON  13.2900 1.5600 13.1350 1.5600 13.1350 1.6800 13.0150 1.6800 13.0150 1.4400
                 13.1700 1.4400 13.1700 1.0600 11.4150 1.0600 11.4150 1.1500 11.2950 1.1500
                 11.2950 0.9100 11.4150 0.9100 11.4150 0.9400 12.9550 0.9400 12.9550 0.7400
                 13.1950 0.7400 13.1950 0.9400 13.2900 0.9400 ;
        POLYGON  12.8050 0.5800 12.4200 0.5800 12.4200 0.8200 11.5350 0.8200 11.5350 0.7900
                 11.1750 0.7900 11.1750 1.2700 11.9050 1.2700 11.9050 1.4400 12.3650 1.4400
                 12.3650 1.5000 12.8050 1.5000 12.8050 1.7400 12.5650 1.7400 12.5650 1.6200
                 12.2450 1.6200 12.2450 1.5600 11.9050 1.5600 11.9050 1.8000 11.7850 1.8000
                 11.7850 1.3900 11.0550 1.3900 11.0550 0.7900 10.9150 0.7900 10.9150 0.9600
                 10.0750 0.9600 10.0750 0.4800 9.4000 0.4800 9.4000 0.5000 9.2650 0.5000 9.2650 1.0550
                 8.8850 1.0550 8.8850 1.1200 8.6450 1.1200 8.6450 1.0000 8.7650 1.0000 8.7650 0.9350
                 9.1450 0.9350 9.1450 0.3800 9.2800 0.3800 9.2800 0.3600 10.1950 0.3600 10.1950 0.8400
                 10.7950 0.8400 10.7950 0.5400 10.9150 0.5400 10.9150 0.6600 11.1750 0.6600
                 11.1750 0.6700 11.6550 0.6700 11.6550 0.7000 12.3000 0.7000 12.3000 0.4600
                 12.8050 0.4600 ;
        POLYGON  12.3850 1.8600 12.2650 1.8600 12.2650 2.0400 11.9100 2.0400 11.9100 2.1100
                 10.9950 2.1100 10.9950 1.9900 10.9750 1.9900 10.9750 1.7500 11.0950 1.7500
                 11.0950 1.8700 11.1150 1.8700 11.1150 1.9900 11.7900 1.9900 11.7900 1.9200
                 12.1450 1.9200 12.1450 1.7400 12.3850 1.7400 ;
        POLYGON  11.5150 1.8700 11.3950 1.8700 11.3950 1.6300 10.6750 1.6300 10.6750 1.8700
                 10.5550 1.8700 10.5550 1.5100 11.5150 1.5100 ;
        POLYGON  10.8750 2.2500 10.3700 2.2500 10.3700 2.1100 9.9250 2.1100 9.9250 2.1300 8.3350 2.1300
                 8.3350 2.1700 3.9750 2.1700 3.9750 1.6900 3.4950 1.6900 3.4950 2.1100 2.3750 2.1100
                 2.3750 2.2500 2.1350 2.2500 2.1350 2.1300 2.1700 2.1300 2.1700 1.8200 1.4950 1.8200
                 1.4950 1.8700 1.3750 1.8700 1.3750 1.8200 1.0250 1.8200 1.0250 1.9600 0.7850 1.9600
                 0.7850 1.8400 0.9050 1.8400 0.9050 1.7000 1.3750 1.7000 1.3750 0.6800 1.6750 0.6800
                 1.6750 0.8000 1.4950 0.8000 1.4950 1.7000 2.2900 1.7000 2.2900 1.9900 3.3750 1.9900
                 3.3750 1.5700 4.0950 1.5700 4.0950 2.0500 8.2150 2.0500 8.2150 2.0100 9.8050 2.0100
                 9.8050 1.9900 10.4900 1.9900 10.4900 2.1300 10.8750 2.1300 ;
        POLYGON  10.4650 1.2500 9.7450 1.2500 9.7450 1.6750 9.7150 1.6750 9.7150 1.8700 9.5950 1.8700
                 9.5950 1.5550 9.6250 1.5550 9.6250 0.6000 9.9550 0.6000 9.9550 0.7200 9.7450 0.7200
                 9.7450 1.1300 10.4650 1.1300 ;
        POLYGON  8.5250 0.4800 7.8750 0.4800 7.8750 0.8200 6.7850 0.8200 6.7850 0.8600 6.5650 0.8600
                 6.5650 1.5700 7.6450 1.5700 7.6450 1.2500 7.8850 1.2500 7.8850 1.3700 7.7650 1.3700
                 7.7650 1.6900 6.4450 1.6900 6.4450 0.7400 6.6650 0.7400 6.6650 0.6200 6.7850 0.6200
                 6.7850 0.7000 7.7550 0.7000 7.7550 0.3600 8.5250 0.3600 ;
        POLYGON  8.4050 1.6900 8.0050 1.6900 8.0050 1.9300 4.7950 1.9300 4.7950 1.6700 4.9150 1.6700
                 4.9150 0.6200 5.0350 0.6200 5.0350 1.8100 7.8850 1.8100 7.8850 1.5700 8.2850 1.5700
                 8.2850 0.8000 8.1450 0.8000 8.1450 0.6800 8.4050 0.6800 ;
        POLYGON  6.3250 1.6900 6.0850 1.6900 6.0850 1.5700 6.1950 1.5700 6.1950 0.9200 5.5950 0.9200
                 5.5950 1.1400 5.4750 1.1400 5.4750 0.8000 6.1950 0.8000 6.1950 0.6800 6.1450 0.6800
                 6.1450 0.4400 6.2650 0.4400 6.2650 0.5600 6.3150 0.5600 6.3150 1.5700 6.3250 1.5700 ;
        POLYGON  5.4250 0.6800 5.3550 0.6800 5.3550 1.5700 5.3950 1.5700 5.3950 1.6900 5.1550 1.6900
                 5.1550 1.5700 5.2350 1.5700 5.2350 0.5000 4.7950 0.5000 4.7950 1.5500 4.6750 1.5500
                 4.6750 0.5000 4.0950 0.5000 4.0950 0.9700 3.3750 0.9700 3.3750 0.5000 2.5350 0.5000
                 2.5350 1.2200 2.5950 1.2200 2.5950 1.3400 2.3550 1.3400 2.3550 1.2200 2.4150 1.2200
                 2.4150 0.3800 2.9350 0.3800 2.9350 0.3600 3.1750 0.3600 3.1750 0.3800 3.4950 0.3800
                 3.4950 0.8500 3.9750 0.8500 3.9750 0.3800 4.1750 0.3800 4.1750 0.3600 4.4150 0.3600
                 4.4150 0.3800 5.4250 0.3800 ;
        POLYGON  4.5550 0.8000 4.4950 0.8000 4.4950 1.8700 4.3750 1.8700 4.3750 1.2100 3.3950 1.2100
                 3.3950 1.0900 4.3750 1.0900 4.3750 0.8000 4.3150 0.8000 4.3150 0.6800 4.5550 0.6800 ;
        POLYGON  4.0750 1.4500 3.2550 1.4500 3.2550 1.8700 3.1350 1.8700 3.1350 0.6200 3.2550 0.6200
                 3.2550 1.3300 4.0750 1.3300 ;
        POLYGON  2.8950 0.8000 2.8350 0.8000 2.8350 1.8700 2.7150 1.8700 2.7150 1.5800 1.7750 1.5800
                 1.7750 1.3100 1.8950 1.3100 1.8950 1.4600 2.7150 1.4600 2.7150 0.8000 2.6550 0.8000
                 2.6550 0.6800 2.8950 0.6800 ;
        POLYGON  1.1050 1.5800 0.9850 1.5800 0.9850 1.1800 0.3750 1.1800 0.3750 1.0600 0.9850 1.0600
                 0.9850 0.6800 1.1050 0.6800 ;
    END
END SEDFFTRXL

MACRO SEDFFTRX4
    CLASS CORE ;
    FOREIGN SEDFFTRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 17.4000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8600 0.3900 1.9800 1.4100 ;
        RECT  0.9000 0.3900 1.9800 0.5100 ;
        RECT  0.3000 0.9700 1.2200 1.0900 ;
        RECT  0.9000 0.3900 1.0200 1.0900 ;
        RECT  0.3050 0.9400 0.5650 1.0900 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2300 0.8800 1.4700 ;
        RECT  0.5950 1.2100 0.8550 1.4700 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1700 1.1750 8.3400 1.4350 ;
        RECT  7.9100 1.3000 8.3400 1.4200 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.0650 1.4700 13.3250 1.7400 ;
        RECT  13.0850 1.3400 13.3250 1.7400 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  15.2750 1.3200 16.2400 1.4400 ;
        RECT  16.1200 1.0600 16.2400 1.4400 ;
        RECT  16.0200 1.1750 16.2400 1.4400 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  16.8650 1.0000 16.9850 1.2400 ;
        RECT  16.6000 1.0000 16.9850 1.1450 ;
        RECT  16.6000 0.8850 16.7500 1.1450 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8200 0.7200 10.0200 0.8400 ;
        RECT  9.4950 1.5200 9.6150 1.8000 ;
        RECT  9.0050 1.5200 9.6150 1.6400 ;
        RECT  8.4750 1.6200 9.2650 1.6700 ;
        RECT  8.4750 1.6200 9.1600 1.7400 ;
        RECT  9.0400 0.7200 9.1600 1.7400 ;
        RECT  8.4750 1.6200 8.7150 1.8000 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7400 0.7200 11.9400 0.8400 ;
        RECT  11.3550 1.6200 11.5950 1.7400 ;
        RECT  10.7450 1.5200 11.4750 1.6400 ;
        RECT  10.3950 1.6200 11.0050 1.6700 ;
        RECT  10.3950 1.6200 10.9800 1.7400 ;
        RECT  10.8600 0.7200 10.9800 1.7400 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 17.4000 0.1800 ;
        RECT  16.6850 -0.1800 16.8050 0.4000 ;
        RECT  15.1150 0.6000 15.3550 0.7200 ;
        RECT  15.1150 -0.1800 15.2350 0.7200 ;
        RECT  14.7850 -0.1800 14.9050 0.4000 ;
        RECT  13.5900 -0.1800 13.8300 0.3800 ;
        RECT  12.1800 -0.1800 12.4200 0.3600 ;
        RECT  11.2200 -0.1800 11.4600 0.3600 ;
        RECT  10.2600 -0.1800 10.5000 0.3600 ;
        RECT  9.3000 -0.1800 9.5400 0.3600 ;
        RECT  8.3400 -0.1800 8.5800 0.3600 ;
        RECT  6.9850 0.5800 7.2250 0.7000 ;
        RECT  6.9850 -0.1800 7.1050 0.7000 ;
        RECT  6.1450 0.5800 6.3850 0.7000 ;
        RECT  6.1450 -0.1800 6.2650 0.7000 ;
        RECT  4.2650 -0.1800 4.5050 0.3200 ;
        RECT  2.1400 -0.1800 2.2600 0.8100 ;
        RECT  0.5600 -0.1800 0.6800 0.8100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 17.4000 2.7900 ;
        RECT  16.6050 2.0800 16.8450 2.2000 ;
        RECT  16.6050 2.0800 16.7250 2.7900 ;
        RECT  13.2650 2.1400 13.3850 2.7900 ;
        RECT  11.8350 2.1600 12.0750 2.2800 ;
        RECT  11.8350 2.1600 11.9550 2.7900 ;
        RECT  10.8750 2.1000 11.1150 2.2200 ;
        RECT  10.8750 2.1000 10.9950 2.7900 ;
        RECT  9.9150 2.1600 10.1550 2.2800 ;
        RECT  9.9150 2.1600 10.0350 2.7900 ;
        RECT  8.9550 2.1600 9.1950 2.2800 ;
        RECT  8.9550 2.1600 9.0750 2.7900 ;
        RECT  7.9950 2.1600 8.2350 2.2800 ;
        RECT  7.9950 2.1600 8.1150 2.7900 ;
        RECT  7.1250 2.2000 7.3650 2.7900 ;
        RECT  6.1850 2.2800 6.4250 2.7900 ;
        RECT  4.0250 2.2200 4.1450 2.7900 ;
        RECT  2.3400 2.2900 2.5800 2.7900 ;
        RECT  0.6200 1.8300 0.8600 1.9500 ;
        RECT  0.6200 1.8300 0.7400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  17.2650 1.8600 16.7350 1.8600 16.7350 1.9600 16.4700 1.9600 16.4700 2.2400
                 15.6150 2.2400 15.6150 2.1200 16.3500 2.1200 16.3500 1.8400 16.6150 1.8400
                 16.6150 1.7400 17.1450 1.7400 17.1450 0.6800 17.2650 0.6800 ;
        POLYGON  16.4800 1.6800 16.1450 1.6800 16.1450 1.5600 16.3600 1.5600 16.3600 0.9200
                 16.2050 0.9200 16.2050 0.4800 15.6050 0.4800 15.6050 0.9600 14.8100 0.9600
                 14.8100 1.1800 14.5700 1.1800 14.5700 1.0600 14.6900 1.0600 14.6900 0.8400
                 15.4850 0.8400 15.4850 0.3600 16.3250 0.3600 16.3250 0.8000 16.4800 0.8000 ;
        POLYGON  15.9950 0.7200 15.8450 0.7200 15.8450 1.2000 15.1550 1.2000 15.1550 1.5600
                 15.9350 1.5600 15.9350 1.8600 15.8150 1.8600 15.8150 1.6800 15.1550 1.6800
                 15.1550 1.8000 14.9150 1.8000 14.9150 1.6800 15.0350 1.6800 15.0350 1.4200
                 13.5650 1.4200 13.5650 1.9800 13.4850 1.9800 13.4850 2.0200 12.9550 2.0200
                 12.9550 2.0400 12.0400 2.0400 12.0400 1.9800 10.3050 1.9800 10.3050 2.0400
                 7.6550 2.0400 7.6550 2.0800 6.0650 2.0800 6.0650 2.2400 4.2650 2.2400 4.2650 2.1000
                 3.9050 2.1000 3.9050 2.1700 2.1400 2.1700 2.1400 2.1500 2.0200 2.1500 2.0200 2.0300
                 2.2600 2.0300 2.2600 2.0500 3.7850 2.0500 3.7850 1.9800 4.3850 1.9800 4.3850 2.1200
                 5.9450 2.1200 5.9450 1.9600 7.5350 1.9600 7.5350 1.9200 10.1850 1.9200 10.1850 1.8600
                 12.1600 1.8600 12.1600 1.9200 12.8350 1.9200 12.8350 1.9000 13.3650 1.9000
                 13.3650 1.8600 13.4450 1.8600 13.4450 1.3000 14.1900 1.3000 14.1900 0.8600
                 14.0700 0.8600 14.0700 0.7400 14.3100 0.7400 14.3100 1.3000 15.0350 1.3000
                 15.0350 1.0800 15.7250 1.0800 15.7250 0.6000 15.9950 0.6000 ;
        POLYGON  15.5750 1.9200 15.4550 1.9200 15.4550 2.0800 14.2250 2.0800 14.2250 1.9000
                 14.1050 1.9000 14.1050 1.7800 14.3450 1.7800 14.3450 1.9600 15.3350 1.9600
                 15.3350 1.8000 15.5750 1.8000 ;
        POLYGON  14.7050 1.8400 14.5850 1.8400 14.5850 1.6600 13.9850 1.6600 13.9850 1.7800
                 13.6850 1.7800 13.6850 1.6600 13.8650 1.6600 13.8650 1.5400 14.7050 1.5400 ;
        POLYGON  14.4500 0.5400 14.0700 0.5400 14.0700 0.6200 13.3500 0.6200 13.3500 0.5600
                 12.9400 0.5600 12.9400 0.6000 12.4100 0.6000 12.4100 1.2400 12.2900 1.2400
                 12.2900 0.6000 8.7000 0.6000 8.7000 0.9800 8.9200 0.9800 8.9200 1.2200 8.5800 1.2200
                 8.5800 1.4600 8.4600 1.4600 8.4600 1.1000 8.5800 1.1000 8.5800 0.6000 7.5400 0.6000
                 7.5400 0.9400 6.7450 0.9400 6.7450 1.3000 6.7650 1.3000 6.7650 1.4800 6.8850 1.4800
                 6.8850 1.6000 6.6450 1.6000 6.6450 1.4200 6.0050 1.4200 6.0050 1.1800 6.1250 1.1800
                 6.1250 1.3000 6.6250 1.3000 6.6250 0.6200 6.7450 0.6200 6.7450 0.8200 7.4200 0.8200
                 7.4200 0.4800 12.8200 0.4800 12.8200 0.4400 13.4700 0.4400 13.4700 0.5000
                 13.9500 0.5000 13.9500 0.4200 14.4500 0.4200 ;
        POLYGON  13.7900 1.1800 12.9450 1.1800 12.9450 1.7800 12.7050 1.7800 12.7050 1.6600
                 12.8250 1.6600 12.8250 0.9600 13.1100 0.9600 13.1100 0.6800 13.2300 0.6800
                 13.2300 1.0600 13.7900 1.0600 ;
        POLYGON  12.9000 0.8400 12.7050 0.8400 12.7050 1.4800 12.4950 1.4800 12.4950 1.8000
                 12.3750 1.8000 12.3750 1.4800 11.6200 1.4800 11.6200 1.2400 11.7400 1.2400
                 11.7400 1.3600 12.5850 1.3600 12.5850 0.7200 12.9000 0.7200 ;
        POLYGON  8.0500 1.1800 7.7900 1.1800 7.7900 1.6800 7.6950 1.6800 7.6950 1.8000 7.1500 1.8000
                 7.1500 1.8400 5.8250 1.8400 5.8250 2.0000 4.5050 2.0000 4.5050 1.6800 3.8450 1.6800
                 3.8450 1.5000 3.7800 1.5000 3.7800 1.2600 3.9000 1.2600 3.9000 1.3800 3.9650 1.3800
                 3.9650 1.5600 4.6250 1.5600 4.6250 1.8800 5.1050 1.8800 5.1050 1.4400 4.9850 1.4400
                 4.9850 1.3200 5.2250 1.3200 5.2250 1.8800 5.7050 1.8800 5.7050 1.1800 5.5850 1.1800
                 5.5850 1.0600 5.8250 1.0600 5.8250 1.7200 7.0300 1.7200 7.0300 1.6800 7.5750 1.6800
                 7.5750 1.5600 7.6700 1.5600 7.6700 1.0600 7.8100 1.0600 7.8100 0.7200 8.0500 0.7200 ;
        POLYGON  6.5050 1.1800 6.3850 1.1800 6.3850 0.9400 5.4650 0.9400 5.4650 1.6400 5.5850 1.6400
                 5.5850 1.7600 5.3450 1.7600 5.3450 0.6200 5.4650 0.6200 5.4650 0.8200 6.5050 0.8200 ;
        POLYGON  5.2250 1.1200 4.9850 1.1200 4.9850 1.0000 5.1050 1.0000 5.1050 0.5600 4.0250 0.5600
                 4.0250 0.5000 3.4200 0.5000 3.4200 1.5000 3.3000 1.5000 3.3000 0.5000 2.8900 0.5000
                 2.8900 0.5700 2.6800 0.5700 2.6800 0.6900 2.7500 0.6900 2.7500 1.5700 2.9400 1.5700
                 2.9400 1.6900 2.6300 1.6900 2.6300 0.8100 2.5600 0.8100 2.5600 0.4500 2.7700 0.4500
                 2.7700 0.3800 3.7050 0.3800 3.7050 0.3600 3.9450 0.3600 3.9450 0.3800 4.1450 0.3800
                 4.1450 0.4400 5.2250 0.4400 ;
        POLYGON  4.9850 0.8000 4.8650 0.8000 4.8650 1.6400 4.9850 1.6400 4.9850 1.7600 4.7450 1.7600
                 4.7450 1.4400 4.0850 1.4400 4.0850 1.3200 4.7450 1.3200 4.7450 0.6800 4.9850 0.6800 ;
        POLYGON  4.6250 1.1200 3.6600 1.1200 3.6600 1.6200 3.7250 1.6200 3.7250 1.8600 3.6050 1.8600
                 3.6050 1.7400 3.5400 1.7400 3.5400 0.6800 3.7800 0.6800 3.7800 0.8000 3.6600 0.8000
                 3.6600 1.0000 4.6250 1.0000 ;
        POLYGON  3.3050 1.9300 2.3900 1.9300 2.3900 1.9100 1.6000 1.9100 1.6000 1.5500 1.6200 1.5500
                 1.6200 0.7500 1.1400 0.7500 1.1400 0.6300 1.7400 0.6300 1.7400 1.6700 1.7200 1.6700
                 1.7200 1.7900 2.5100 1.7900 2.5100 1.8100 3.0600 1.8100 3.0600 0.6200 3.1800 0.6200
                 3.1800 1.6200 3.3050 1.6200 ;
        POLYGON  1.5000 1.4300 1.4800 1.4300 1.4800 1.7100 0.3200 1.7100 0.3200 1.8300 0.2000 1.8300
                 0.2000 1.7100 0.0600 1.7100 0.0600 0.6900 0.1400 0.6900 0.1400 0.5700 0.2600 0.5700
                 0.2600 0.8100 0.1800 0.8100 0.1800 1.5900 1.3600 1.5900 1.3600 1.3100 1.3800 1.3100
                 1.3800 1.1900 1.5000 1.1900 ;
    END
END SEDFFTRX4

MACRO SEDFFTRX2
    CLASS CORE ;
    FOREIGN SEDFFTRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.7900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8600 0.3900 1.9800 1.4100 ;
        RECT  0.9000 0.3900 1.9800 0.5100 ;
        RECT  0.3000 0.9700 1.2200 1.0900 ;
        RECT  0.9000 0.3900 1.0200 1.0900 ;
        RECT  0.3050 0.9400 0.5650 1.0900 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2300 0.8800 1.4700 ;
        RECT  0.5950 1.2100 0.8550 1.4700 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3200 1.1750 7.4700 1.5850 ;
        RECT  7.3500 1.1000 7.4700 1.5850 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.2300 10.7350 1.4800 ;
        RECT  10.4550 1.2300 10.7150 1.5000 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.7450 1.1800 13.8650 1.4200 ;
        RECT  12.7500 1.2600 13.8650 1.3800 ;
        RECT  13.3550 1.2300 13.6150 1.3800 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  14.2250 1.1500 14.4850 1.4200 ;
        RECT  14.2250 1.0200 14.4650 1.4200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0900 1.1750 8.3400 1.4350 ;
        RECT  8.0700 0.7400 8.3100 0.8600 ;
        RECT  8.0900 0.7400 8.2100 1.4800 ;
        RECT  8.0400 1.3600 8.1600 1.6800 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0000 0.7400 9.2700 0.8600 ;
        RECT  9.0000 0.7400 9.1200 1.6800 ;
        RECT  8.7700 1.1750 9.1200 1.4350 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.7900 0.1800 ;
        RECT  14.1150 -0.1800 14.2350 0.8200 ;
        RECT  12.4300 0.5100 12.6700 0.6300 ;
        RECT  12.4300 -0.1800 12.5500 0.6300 ;
        RECT  12.1000 -0.1800 12.2200 0.6300 ;
        RECT  10.8600 -0.1800 11.1000 0.3200 ;
        RECT  9.5100 -0.1800 9.7500 0.3800 ;
        RECT  8.5500 -0.1800 8.7900 0.3800 ;
        RECT  7.5900 -0.1800 7.8300 0.3400 ;
        RECT  6.2400 0.5300 6.4800 0.6500 ;
        RECT  6.2400 -0.1800 6.3600 0.6500 ;
        RECT  4.2400 0.5500 4.4800 0.6700 ;
        RECT  4.3600 -0.1800 4.4800 0.6700 ;
        RECT  2.1400 -0.1800 2.2600 0.8100 ;
        RECT  0.5600 -0.1800 0.6800 0.8100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.7900 2.7900 ;
        RECT  14.0550 2.1600 14.1750 2.7900 ;
        RECT  10.8750 2.0100 10.9950 2.7900 ;
        RECT  10.7550 2.0100 10.9950 2.1300 ;
        RECT  9.4800 2.0800 9.6000 2.7900 ;
        RECT  8.4600 2.0400 8.7000 2.1600 ;
        RECT  8.4600 2.0400 8.5800 2.7900 ;
        RECT  7.5600 2.2100 7.6800 2.7900 ;
        RECT  6.1700 2.2900 6.4100 2.7900 ;
        RECT  4.0100 2.2300 4.1300 2.7900 ;
        RECT  2.3400 2.2900 2.5800 2.7900 ;
        RECT  0.6200 1.8300 0.8600 1.9500 ;
        RECT  0.6200 1.8300 0.7400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.7250 1.6600 14.6550 1.6600 14.6550 1.9000 14.1400 1.9000 14.1400 2.0400
                 13.6100 2.0400 13.6100 2.1800 13.1050 2.1800 13.1050 2.0600 13.4900 2.0600
                 13.4900 1.9200 14.0200 1.9200 14.0200 1.7800 14.5350 1.7800 14.5350 1.5400
                 14.6050 1.5400 14.6050 0.9000 14.5350 0.9000 14.5350 0.5800 14.6550 0.5800
                 14.6550 0.7800 14.7250 0.7800 ;
        POLYGON  14.1050 1.6600 13.8150 1.6600 13.8150 1.7800 13.6950 1.7800 13.6950 1.5400
                 13.9850 1.5400 13.9850 1.0600 13.6950 1.0600 13.6950 0.4800 12.9100 0.4800
                 12.9100 0.8700 12.0350 0.8700 12.0350 1.2600 11.9150 1.2600 11.9150 0.7500
                 12.7900 0.7500 12.7900 0.3600 13.8150 0.3600 13.8150 0.9400 14.1050 0.9400 ;
        POLYGON  13.4250 1.8000 13.3050 1.8000 13.3050 1.6200 12.6300 1.6200 12.6300 1.6800
                 12.5850 1.6800 12.5850 1.8000 12.4650 1.8000 12.4650 1.5000 10.9750 1.5000
                 10.9750 1.8900 10.6350 1.8900 10.6350 2.2500 9.7200 2.2500 9.7200 1.9200 7.4550 1.9200
                 7.4550 2.0900 6.0500 2.0900 6.0500 2.2500 4.2500 2.2500 4.2500 2.1100 3.8900 2.1100
                 3.8900 2.1700 2.1400 2.1700 2.1400 2.1500 2.0200 2.1500 2.0200 2.0300 2.2600 2.0300
                 2.2600 2.0500 3.7700 2.0500 3.7700 1.9900 4.3700 1.9900 4.3700 2.1300 5.9300 2.1300
                 5.9300 1.9700 7.3350 1.9700 7.3350 1.8000 9.8400 1.8000 9.8400 2.1300 10.5150 2.1300
                 10.5150 1.7700 10.8550 1.7700 10.8550 1.3800 11.4600 1.3800 11.4600 0.8600
                 11.3400 0.8600 11.3400 0.7400 11.5800 0.7400 11.5800 1.3800 12.5100 1.3800
                 12.5100 0.9900 13.1300 0.9900 13.1300 0.6000 13.3700 0.6000 13.3700 0.7200
                 13.2500 0.7200 13.2500 1.1100 12.6300 1.1100 12.6300 1.5000 13.4250 1.5000 ;
        POLYGON  13.0650 1.8600 12.9450 1.8600 12.9450 2.0400 12.5700 2.0400 12.5700 2.2500
                 11.6550 2.2500 11.6550 1.9500 11.7750 1.9500 11.7750 2.1300 12.4500 2.1300
                 12.4500 1.9200 12.8250 1.9200 12.8250 1.7400 13.0650 1.7400 ;
        POLYGON  12.2550 2.0100 12.0150 2.0100 12.0150 1.8300 11.5350 1.8300 11.5350 2.0100
                 11.1750 2.0100 11.1750 1.8900 11.4150 1.8900 11.4150 1.7100 12.1350 1.7100
                 12.1350 1.8900 12.2550 1.8900 ;
        POLYGON  11.7400 0.5200 11.3950 0.5200 11.3950 0.5600 10.0700 0.5600 10.0700 0.6200
                 7.9500 0.6200 7.9500 0.9800 7.9700 0.9800 7.9700 1.2400 7.8500 1.2400 7.8500 1.1000
                 7.8300 1.1000 7.8300 0.6200 6.9000 0.6200 6.9000 0.8600 6.7900 0.8600 6.7900 1.4900
                 6.8700 1.4900 6.8700 1.6100 6.6300 1.6100 6.6300 1.4500 5.9300 1.4500 5.9300 1.3300
                 6.6700 1.3300 6.6700 0.7400 6.7800 0.7400 6.7800 0.5000 9.8700 0.5000 9.8700 0.4000
                 10.1100 0.4000 10.1100 0.4400 11.2750 0.4400 11.2750 0.4000 11.7400 0.4000 ;
        POLYGON  11.1350 1.1800 10.8550 1.1800 10.8550 1.1100 10.3350 1.1100 10.3350 1.8900
                 10.3950 1.8900 10.3950 2.0100 10.1550 2.0100 10.1550 1.8900 10.2150 1.8900
                 10.2150 0.9800 10.4400 0.9800 10.4400 0.6800 10.5600 0.6800 10.5600 0.9900
                 10.9750 0.9900 10.9750 1.0600 11.1350 1.0600 ;
        POLYGON  10.2300 0.8600 10.0950 0.8600 10.0950 1.3000 10.0250 1.3000 10.0250 1.6800
                 9.9050 1.6800 9.9050 1.3000 9.2400 1.3000 9.2400 1.1800 9.9750 1.1800 9.9750 0.7400
                 10.2300 0.7400 ;
        POLYGON  7.3500 0.8600 7.2000 0.8600 7.2000 1.8500 5.8100 1.8500 5.8100 2.0100 4.4900 2.0100
                 4.4900 1.6900 3.8100 1.6900 3.8100 1.2700 3.9300 1.2700 3.9300 1.5700 4.6100 1.5700
                 4.6100 1.8900 5.0900 1.8900 5.0900 1.4500 5.0700 1.4500 5.0700 1.3300 5.3100 1.3300
                 5.3100 1.4500 5.2100 1.4500 5.2100 1.8900 5.6900 1.8900 5.6900 1.1300 5.6800 1.1300
                 5.6800 1.0100 5.9200 1.0100 5.9200 1.1300 5.8100 1.1300 5.8100 1.7300 7.0800 1.7300
                 7.0800 0.7400 7.3500 0.7400 ;
        POLYGON  6.5500 1.2000 6.4300 1.2000 6.4300 0.8900 5.5600 0.8900 5.5600 1.6500 5.5700 1.6500
                 5.5700 1.7700 5.3300 1.7700 5.3300 1.6500 5.4400 1.6500 5.4400 0.7400 5.4800 0.7400
                 5.4800 0.6200 5.6000 0.6200 5.6000 0.7400 5.7550 0.7400 5.7550 0.7700 6.5500 0.7700 ;
        POLYGON  5.3200 1.1800 5.2000 1.1800 5.2000 0.5600 4.7200 0.5600 4.7200 0.9100 4.0000 0.9100
                 4.0000 0.5000 3.4200 0.5000 3.4200 1.5100 3.3000 1.5100 3.3000 0.5000 2.8900 0.5000
                 2.8900 0.5700 2.6800 0.5700 2.6800 0.6900 2.7400 0.6900 2.7400 1.5700 2.9400 1.5700
                 2.9400 1.6900 2.6200 1.6900 2.6200 0.8100 2.5600 0.8100 2.5600 0.4500 2.7700 0.4500
                 2.7700 0.3800 3.6800 0.3800 3.6800 0.3600 3.9200 0.3600 3.9200 0.3800 4.1200 0.3800
                 4.1200 0.7900 4.6000 0.7900 4.6000 0.4400 5.3200 0.4400 ;
        POLYGON  5.0800 1.1500 4.9500 1.1500 4.9500 1.6500 4.9700 1.6500 4.9700 1.7700 4.7300 1.7700
                 4.7300 1.6500 4.8300 1.6500 4.8300 1.4500 4.1100 1.4500 4.1100 1.3300 4.8300 1.3300
                 4.8300 1.0300 4.8400 1.0300 4.8400 0.6800 5.0800 0.6800 ;
        POLYGON  4.7100 1.1500 3.6900 1.1500 3.6900 1.8300 3.5700 1.8300 3.5700 0.8000 3.5400 0.8000
                 3.5400 0.6800 3.7800 0.6800 3.7800 0.8000 3.6900 0.8000 3.6900 1.0300 4.7100 1.0300 ;
        POLYGON  3.2700 1.9300 2.3800 1.9300 2.3800 1.9100 1.6000 1.9100 1.6000 1.5500 1.6200 1.5500
                 1.6200 0.7500 1.1400 0.7500 1.1400 0.6300 1.7400 0.6300 1.7400 1.6700 1.7200 1.6700
                 1.7200 1.7900 2.5000 1.7900 2.5000 1.8100 3.0600 1.8100 3.0600 0.6200 3.1800 0.6200
                 3.1800 1.6300 3.2700 1.6300 ;
        POLYGON  1.5000 1.4300 1.4800 1.4300 1.4800 1.7100 0.3200 1.7100 0.3200 1.8300 0.2000 1.8300
                 0.2000 1.7100 0.0600 1.7100 0.0600 0.6900 0.1400 0.6900 0.1400 0.5700 0.2600 0.5700
                 0.2600 0.8100 0.1800 0.8100 0.1800 1.5900 1.3600 1.5900 1.3600 1.3100 1.3800 1.3100
                 1.3800 1.1900 1.5000 1.1900 ;
    END
END SEDFFTRX2

MACRO SEDFFTRX1
    CLASS CORE ;
    FOREIGN SEDFFTRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.7900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8700 1.1300 6.1000 1.4400 ;
        END
    END CK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2000 0.8100 8.3200 1.2000 ;
        RECT  7.1150 0.8100 8.3200 0.9300 ;
        RECT  7.1150 0.8100 7.2350 1.2000 ;
        RECT  6.9750 0.9400 7.2350 1.0900 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5600 1.0500 7.7600 1.4350 ;
        RECT  7.5600 1.0500 7.6800 1.4500 ;
        END
    END SI
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.2100 1.3500 10.4500 1.5050 ;
        RECT  10.2200 1.3500 10.3700 1.7250 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.4100 1.4650 13.5600 1.7250 ;
        RECT  13.4100 1.2700 13.5300 1.7250 ;
        RECT  12.4700 1.2700 13.5300 1.3900 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  14.2400 1.0400 14.3600 1.2800 ;
        RECT  14.0200 1.1600 14.3600 1.2800 ;
        RECT  13.9900 1.1750 14.1400 1.4350 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6200 1.1750 9.7900 1.4350 ;
        RECT  9.4000 1.4900 9.7400 1.6100 ;
        RECT  9.6200 0.6800 9.7400 1.6100 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.7900 0.1800 ;
        RECT  14.1000 -0.1800 14.2200 0.9200 ;
        RECT  12.2100 0.5500 12.4500 0.6700 ;
        RECT  12.2100 -0.1800 12.3300 0.6700 ;
        RECT  11.6700 0.5500 11.9100 0.6700 ;
        RECT  11.6700 -0.1800 11.7900 0.6700 ;
        RECT  10.5500 0.6000 10.7900 0.7200 ;
        RECT  10.6700 -0.1800 10.7900 0.7200 ;
        RECT  9.1400 -0.1800 9.2600 0.7300 ;
        RECT  7.2800 0.3300 7.5200 0.4500 ;
        RECT  7.2800 -0.1800 7.4000 0.4500 ;
        RECT  5.8000 -0.1800 5.9200 0.7700 ;
        RECT  3.6900 0.6100 3.9300 0.7300 ;
        RECT  3.8100 -0.1800 3.9300 0.7300 ;
        RECT  1.9900 -0.1800 2.1100 0.8600 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.7900 2.7900 ;
        RECT  14.1600 2.0000 14.2800 2.7900 ;
        RECT  10.4000 2.2300 10.6400 2.7900 ;
        RECT  8.9200 1.9700 9.1600 2.0900 ;
        RECT  8.9200 1.9700 9.0400 2.7900 ;
        RECT  7.2800 2.2900 7.5200 2.7900 ;
        RECT  5.8000 2.2900 6.0400 2.7900 ;
        RECT  3.8700 1.8100 3.9900 2.7900 ;
        RECT  3.7500 1.8100 3.9900 1.9300 ;
        RECT  1.8500 1.9400 2.0900 2.0600 ;
        RECT  1.8500 1.9400 1.9700 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.6550 1.8400 13.8600 1.8400 13.8600 2.0500 13.0500 2.0500 13.0500 2.1900
                 12.8100 2.1900 12.8100 2.0700 12.9300 2.0700 12.9300 1.9300 13.7400 1.9300
                 13.7400 1.7200 14.5350 1.7200 14.5350 0.9200 14.5200 0.9200 14.5200 0.6800
                 14.6400 0.6800 14.6400 0.8000 14.6550 0.8000 ;
        POLYGON  13.8000 1.6000 13.6800 1.6000 13.6800 1.1500 11.5600 1.1500 11.5600 1.0300
                 13.6800 1.0300 13.6800 0.6800 13.8000 0.6800 ;
        POLYGON  13.1300 1.8100 13.0100 1.8100 13.0100 1.6300 12.2900 1.6300 12.2900 1.8100
                 12.1700 1.8100 12.1700 1.3900 11.3200 1.3900 11.3200 0.9100 11.1500 0.9100
                 11.1500 0.9600 10.3100 0.9600 10.3100 0.4800 9.6350 0.4800 9.6350 0.5600 9.5000 0.5600
                 9.5000 0.9700 9.0400 0.9700 9.0400 1.2000 8.9200 1.2000 8.9200 0.8500 9.3800 0.8500
                 9.3800 0.4400 9.5150 0.4400 9.5150 0.3600 10.4300 0.3600 10.4300 0.8400 11.0300 0.8400
                 11.0300 0.5400 11.1500 0.5400 11.1500 0.6600 11.4400 0.6600 11.4400 0.7900
                 12.5850 0.7900 12.5850 0.5500 13.0900 0.5500 13.0900 0.6700 12.7050 0.6700
                 12.7050 0.9100 11.4400 0.9100 11.4400 1.2700 12.2900 1.2700 12.2900 1.5100
                 13.1300 1.5100 ;
        POLYGON  12.7700 1.8700 12.6500 1.8700 12.6500 2.0500 12.1400 2.0500 12.1400 2.1100
                 11.3800 2.1100 11.3800 1.9900 11.3600 1.9900 11.3600 1.7500 11.4800 1.7500
                 11.4800 1.8700 11.5000 1.8700 11.5000 1.9900 12.0200 1.9900 12.0200 1.9300
                 12.5300 1.9300 12.5300 1.7500 12.7700 1.7500 ;
        POLYGON  11.9000 1.8700 11.7800 1.8700 11.7800 1.6300 11.0600 1.6300 11.0600 1.8700
                 10.9400 1.8700 10.9400 1.5100 11.9000 1.5100 ;
        POLYGON  11.2600 2.2500 11.0150 2.2500 11.0150 2.1100 9.6900 2.1100 9.6900 1.8500 8.8000 1.8500
                 8.8000 2.1700 4.1750 2.1700 4.1750 1.6900 3.6300 1.6900 3.6300 2.1100 2.4500 2.1100
                 2.4500 2.2500 2.2100 2.2500 2.2100 2.1300 2.2250 2.1300 2.2250 1.8200 1.5500 1.8200
                 1.5500 1.8700 1.4300 1.8700 1.4300 1.8200 1.0750 1.8200 1.0750 1.9600 0.8350 1.9600
                 0.8350 1.8400 0.9550 1.8400 0.9550 1.7000 1.4300 1.7000 1.4300 1.6300 1.5700 1.6300
                 1.5700 0.6200 1.6900 0.6200 1.6900 1.7000 2.3450 1.7000 2.3450 1.9900 3.5100 1.9900
                 3.5100 1.5700 4.2950 1.5700 4.2950 2.0500 8.6800 2.0500 8.6800 1.7300 9.1600 1.7300
                 9.1600 1.2100 9.2400 1.2100 9.2400 1.0900 9.3600 1.0900 9.3600 1.3300 9.2800 1.3300
                 9.2800 1.7300 9.8100 1.7300 9.8100 1.9900 11.1350 1.9900 11.1350 2.1300 11.2600 2.1300 ;
        POLYGON  10.8400 1.2300 10.0900 1.2300 10.0900 1.6250 10.1000 1.6250 10.1000 1.8700
                 9.9800 1.8700 9.9800 1.7450 9.9700 1.7450 9.9700 0.7200 9.9500 0.7200 9.9500 0.6000
                 10.1900 0.6000 10.1900 0.7200 10.0900 0.7200 10.0900 1.1100 10.8400 1.1100 ;
        POLYGON  8.7600 0.4800 7.7600 0.4800 7.7600 0.6900 6.8550 0.6900 6.8550 1.5700 7.8800 1.5700
                 7.8800 1.1700 8.0000 1.1700 8.0000 1.6900 6.7350 1.6900 6.7350 0.5700 7.6400 0.5700
                 7.6400 0.3600 8.7600 0.3600 ;
        POLYGON  8.5600 1.6900 8.2400 1.6900 8.2400 1.9300 4.9900 1.9300 4.9900 0.8600 4.9300 0.8600
                 4.9300 0.6200 5.0500 0.6200 5.0500 0.7400 5.1100 0.7400 5.1100 1.8100 8.1200 1.8100
                 8.1200 1.5700 8.4400 1.5700 8.4400 0.6200 8.5600 0.6200 ;
        POLYGON  6.4600 1.6900 6.3400 1.6900 6.3400 1.5700 6.2200 1.5700 6.2200 1.0100 5.7500 1.0100
                 5.7500 1.1400 5.6300 1.1400 5.6300 0.8900 6.2200 0.8900 6.2200 0.5300 6.3400 0.5300
                 6.3400 1.4500 6.4600 1.4500 ;
        POLYGON  5.5000 1.6900 5.3800 1.6900 5.3800 0.5300 5.1700 0.5300 5.1700 0.5000 4.8100 0.5000
                 4.8100 1.3100 4.8700 1.3100 4.8700 1.5500 4.7500 1.5500 4.7500 1.4300 4.6900 1.4300
                 4.6900 0.5000 4.1700 0.5000 4.1700 0.9700 3.4500 0.9700 3.4500 0.5000 2.6100 0.5000
                 2.6100 1.2200 2.6700 1.2200 2.6700 1.3400 2.4300 1.3400 2.4300 1.2200 2.4900 1.2200
                 2.4900 0.3800 3.0100 0.3800 3.0100 0.3600 3.2500 0.3600 3.2500 0.3800 3.5700 0.3800
                 3.5700 0.8500 4.0500 0.8500 4.0500 0.3800 4.2500 0.3800 4.2500 0.3600 4.4900 0.3600
                 4.4900 0.3800 5.2900 0.3800 5.2900 0.4100 5.5000 0.4100 ;
        POLYGON  4.5700 1.8700 4.4500 1.8700 4.4500 1.2100 3.4700 1.2100 3.4700 1.0900 4.4500 1.0900
                 4.4500 0.6200 4.5700 0.6200 ;
        POLYGON  4.1500 1.4500 3.3300 1.4500 3.3300 1.8700 3.2100 1.8700 3.2100 0.6200 3.3300 0.6200
                 3.3300 1.3300 4.1500 1.3300 ;
        POLYGON  2.9700 0.8000 2.9100 0.8000 2.9100 1.8700 2.7900 1.8700 2.7900 1.5800 1.8500 1.5800
                 1.8500 1.3100 1.9700 1.3100 1.9700 1.4600 2.7900 1.4600 2.7900 0.8000 2.7300 0.8000
                 2.7300 0.6800 2.9700 0.6800 ;
        POLYGON  1.1550 1.5800 1.0350 1.5800 1.0350 1.1800 0.3750 1.1800 0.3750 1.0600 1.0350 1.0600
                 1.0350 0.6800 1.1550 0.6800 ;
    END
END SEDFFTRX1

MACRO SEDFFHQX8
    CLASS CORE ;
    FOREIGN SEDFFHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.7900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 1.4650 2.7750 2.2100 ;
        RECT  2.6550 0.6800 2.7750 1.0050 ;
        RECT  2.6350 0.8850 2.7550 1.5850 ;
        RECT  0.0700 1.0050 2.7550 1.1250 ;
        RECT  1.8150 0.6800 1.9350 2.2100 ;
        RECT  0.9750 0.6800 1.0950 2.2050 ;
        RECT  0.1350 0.6800 0.2550 2.2050 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 1.1500 5.1500 1.4700 ;
        RECT  4.9100 1.1500 5.1500 1.4650 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.3050 1.2200 10.6650 1.3500 ;
        RECT  10.1650 1.2300 10.4250 1.3950 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.2500 1.1400 12.4000 1.6100 ;
        RECT  12.2550 1.1400 12.3750 1.6400 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.9350 1.2100 14.1950 1.4650 ;
        RECT  13.8550 1.2100 14.1950 1.4400 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  14.3150 0.9700 14.4350 1.2100 ;
        RECT  13.1350 0.9700 14.4350 1.0900 ;
        RECT  13.6150 0.9400 13.9050 1.0900 ;
        RECT  13.6150 0.9200 13.7350 1.1600 ;
        RECT  13.1350 0.9700 13.2550 1.2600 ;
        RECT  13.0550 1.1400 13.1750 1.4400 ;
        END
    END E
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.7900 0.1800 ;
        RECT  14.1150 -0.1800 14.2350 0.8200 ;
        RECT  12.5350 0.6000 12.7750 0.7200 ;
        RECT  12.5350 -0.1800 12.6550 0.7200 ;
        RECT  10.4650 -0.1800 10.5850 0.6500 ;
        RECT  9.5050 -0.1800 9.6250 0.6300 ;
        RECT  7.0700 0.5000 7.3100 0.6200 ;
        RECT  7.0700 -0.1800 7.1900 0.6200 ;
        RECT  5.3700 0.4300 5.6100 0.5500 ;
        RECT  5.4900 -0.1800 5.6100 0.5500 ;
        RECT  3.9150 -0.1800 4.0350 0.6700 ;
        RECT  3.0750 -0.1800 3.1950 0.6700 ;
        RECT  2.2350 -0.1800 2.3550 0.6700 ;
        RECT  1.3950 -0.1800 1.5150 0.6700 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.7900 2.7900 ;
        RECT  13.9350 1.8250 14.0550 2.7900 ;
        RECT  12.4550 2.2800 12.6950 2.7900 ;
        RECT  10.3450 1.9400 10.5850 2.0900 ;
        RECT  10.3450 1.9400 10.4650 2.7900 ;
        RECT  9.5050 2.1400 9.6250 2.7900 ;
        RECT  7.4300 1.9400 7.6700 2.0600 ;
        RECT  7.4300 1.9400 7.5500 2.7900 ;
        RECT  5.0700 2.1100 5.1900 2.7900 ;
        RECT  3.9150 1.5600 4.0350 2.7900 ;
        RECT  3.0750 1.5600 3.1950 2.7900 ;
        RECT  2.2350 1.4650 2.3550 2.7900 ;
        RECT  1.3950 1.4650 1.5150 2.7900 ;
        RECT  0.5550 1.4650 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.6750 1.7050 14.5350 1.7050 14.5350 1.8250 14.4150 1.8250 14.4150 1.7050
                 13.6150 1.7050 13.6150 1.4200 13.3750 1.4200 13.3750 1.3000 13.7350 1.3000
                 13.7350 1.5850 14.5550 1.5850 14.5550 0.8500 14.5350 0.8500 14.5350 0.5800
                 14.6550 0.5800 14.6550 0.7300 14.6750 0.7300 ;
        POLYGON  13.5950 0.8000 13.0150 0.8000 13.0150 1.0200 12.9350 1.0200 12.9350 1.5600
                 13.3350 1.5600 13.3350 2.2100 13.2150 2.2100 13.2150 1.6800 12.8150 1.6800
                 12.8150 1.0200 12.0050 1.0200 12.0050 1.4400 11.8550 1.4400 11.8550 1.6800
                 11.5850 1.6800 11.5850 1.5600 11.7350 1.5600 11.7350 1.3200 11.8850 1.3200
                 11.8850 0.8400 11.7850 0.8400 11.7850 0.6000 11.9050 0.6000 11.9050 0.7200
                 12.0050 0.7200 12.0050 0.9000 12.8950 0.9000 12.8950 0.6800 13.4750 0.6800
                 13.4750 0.5600 13.5950 0.5600 ;
        POLYGON  12.6950 2.1200 12.4300 2.1200 12.4300 2.1600 12.1650 2.1600 12.1650 2.2500
                 10.7200 2.2500 10.7200 1.8200 10.1050 1.8200 10.1050 2.1500 9.9850 2.1500
                 9.9850 1.6350 9.9250 1.6350 9.9250 0.9900 9.9850 0.9900 9.9850 0.6000 10.1050 0.6000
                 10.1050 1.1100 10.0450 1.1100 10.0450 1.5150 10.1050 1.5150 10.1050 1.7000
                 10.8400 1.7000 10.8400 2.1300 12.0450 2.1300 12.0450 2.0400 12.3100 2.0400
                 12.3100 2.0000 12.5750 2.0000 12.5750 1.2200 12.6950 1.2200 ;
        POLYGON  12.2950 0.7800 12.1750 0.7800 12.1750 0.4800 11.6150 0.4800 11.6150 0.9600
                 11.7650 0.9600 11.7650 1.2000 11.6150 1.2000 11.6150 1.3400 11.4650 1.3400
                 11.4650 1.8000 11.9750 1.8000 11.9750 1.7600 12.2150 1.7600 12.2150 1.8800
                 12.0950 1.8800 12.0950 1.9200 11.3450 1.9200 11.3450 1.3400 11.0250 1.3400
                 11.0250 1.2200 11.4950 1.2200 11.4950 0.3600 12.2950 0.3600 ;
        POLYGON  11.3750 0.8900 10.9050 0.8900 10.9050 1.4600 11.1050 1.4600 11.1050 1.5600
                 11.2250 1.5600 11.2250 2.0100 10.9850 2.0100 10.9850 1.5800 10.7850 1.5800
                 10.7850 0.8900 10.2250 0.8900 10.2250 0.4800 9.8650 0.4800 9.8650 0.8700 9.2650 0.8700
                 9.2650 0.5400 8.3100 0.5400 8.3100 0.9100 8.8700 0.9100 8.8700 1.7700 8.7500 1.7700
                 8.7500 1.0300 8.1900 1.0300 8.1900 0.4200 9.3850 0.4200 9.3850 0.7500 9.7450 0.7500
                 9.7450 0.3600 10.3450 0.3600 10.3450 0.7700 11.2550 0.7700 11.2550 0.6000
                 11.3750 0.6000 ;
        POLYGON  9.8050 1.5200 9.6500 1.5200 9.6500 2.0200 9.3850 2.0200 9.3850 2.2500 7.7900 2.2500
                 7.7900 1.8200 7.3100 1.8200 7.3100 2.2500 5.3350 2.2500 5.3350 1.9900 4.4550 1.9900
                 4.4550 2.2100 4.3350 2.2100 4.3350 1.4400 3.6150 1.4400 3.6150 2.2100 3.4950 2.2100
                 3.4950 1.2450 2.8750 1.2450 2.8750 1.1250 3.4950 1.1250 3.4950 0.6200 3.6150 0.6200
                 3.6150 1.3200 4.3950 1.3200 4.3950 0.6200 4.5150 0.6200 4.5150 1.4400 4.4550 1.4400
                 4.4550 1.8700 5.2700 1.8700 5.2700 1.1500 5.3900 1.1500 5.3900 1.8700 5.4550 1.8700
                 5.4550 2.1300 7.1900 2.1300 7.1900 1.7000 7.9100 1.7000 7.9100 2.1300 9.2650 2.1300
                 9.2650 1.9000 9.5300 1.9000 9.5300 1.4000 9.6850 1.4000 9.6850 1.1600 9.8050 1.1600 ;
        POLYGON  9.2600 1.7800 9.1450 1.7800 9.1450 2.0100 8.0300 2.0100 8.0300 1.5800 7.0700 1.5800
                 7.0700 2.0100 5.6300 2.0100 5.6300 1.1500 5.7500 1.1500 5.7500 1.8900 6.4700 1.8900
                 6.4700 0.8600 6.5900 0.8600 6.5900 1.8900 6.9500 1.8900 6.9500 1.4600 7.7100 1.4600
                 7.7100 1.1000 7.5900 1.1000 7.5900 0.9800 7.8300 0.9800 7.8300 1.4600 8.1500 1.4600
                 8.1500 1.8900 8.5100 1.8900 8.5100 1.1500 8.6300 1.1500 8.6300 1.8900 9.0250 1.8900
                 9.0250 0.7800 8.9050 0.7800 8.9050 0.6600 9.1450 0.6600 9.1450 1.5000 9.2600 1.5000 ;
        POLYGON  8.3900 1.7700 8.2700 1.7700 8.2700 1.3400 7.9500 1.3400 7.9500 0.7800 7.5500 0.7800
                 7.5500 0.8600 7.0700 0.8600 7.0700 1.1000 6.9500 1.1000 6.9500 0.7400 7.4300 0.7400
                 7.4300 0.6600 7.7700 0.6600 7.7700 0.5400 7.8900 0.5400 7.8900 0.6600 8.0700 0.6600
                 8.0700 1.2200 8.3900 1.2200 ;
        POLYGON  7.4700 1.3100 7.3500 1.3100 7.3500 1.3400 6.8300 1.3400 6.8300 1.7700 6.7100 1.7700
                 6.7100 0.5400 6.8300 0.5400 6.8300 1.2200 7.2300 1.2200 7.2300 1.1900 7.4700 1.1900 ;
        POLYGON  6.3500 1.7700 6.2300 1.7700 6.2300 0.7800 6.0450 0.7800 6.0450 0.7900 5.1300 0.7900
                 5.1300 0.4800 4.2750 0.4800 4.2750 1.2000 4.1550 1.2000 4.1550 0.3600 5.2500 0.3600
                 5.2500 0.6700 5.9250 0.6700 5.9250 0.6600 6.2300 0.6600 6.2300 0.5400 6.3500 0.5400 ;
        POLYGON  6.1100 1.1500 5.9900 1.1500 5.9900 1.0300 4.7900 1.0300 4.7900 1.5900 4.7650 1.5900
                 4.7650 1.7100 4.6450 1.7100 4.6450 1.4700 4.6700 1.4700 4.6700 0.6000 5.0100 0.6000
                 5.0100 0.7200 4.7900 0.7200 4.7900 0.9100 6.1100 0.9100 ;
    END
END SEDFFHQX8

MACRO SEDFFHQX4
    CLASS CORE ;
    FOREIGN SEDFFHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.6300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 0.6300 1.5150 1.9900 ;
        RECT  0.5550 1.0250 1.5150 1.1450 ;
        RECT  0.5550 0.8850 0.8000 1.1450 ;
        RECT  0.5550 0.6300 0.6750 1.9900 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2750 1.0300 8.3950 1.4400 ;
        RECT  8.1350 1.1500 8.3950 1.3800 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7700 1.1400 9.0050 1.4600 ;
        RECT  8.7700 1.1350 8.9200 1.4600 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7450 1.1800 11.0050 1.4100 ;
        RECT  10.8450 1.0000 10.9650 1.4100 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.4850 1.2100 12.8650 1.4000 ;
        RECT  12.4850 1.2100 12.7450 1.4250 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.0050 0.9700 13.1250 1.2100 ;
        RECT  12.7750 0.9400 13.0350 1.0900 ;
        RECT  11.8450 0.9700 13.1250 1.0900 ;
        RECT  11.7250 1.2800 11.9650 1.4000 ;
        RECT  11.8450 0.9700 11.9650 1.4000 ;
        END
    END E
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.6300 0.1800 ;
        RECT  12.8450 -0.1800 12.9650 0.8200 ;
        RECT  11.2450 -0.1800 11.3650 0.6400 ;
        RECT  8.5250 0.5100 8.7650 0.6300 ;
        RECT  8.5250 -0.1800 8.6450 0.6300 ;
        RECT  7.0700 -0.1800 7.1900 0.7300 ;
        RECT  4.6550 0.4900 4.8950 0.6100 ;
        RECT  4.7750 -0.1800 4.8950 0.6100 ;
        RECT  2.7750 -0.1800 2.8950 0.6800 ;
        RECT  1.8150 -0.1800 1.9350 0.6800 ;
        RECT  0.9750 -0.1800 1.0950 0.6800 ;
        RECT  0.1350 -0.1800 0.2550 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.6300 2.7900 ;
        RECT  12.6850 1.7850 12.8050 2.7900 ;
        RECT  11.3050 1.7700 11.4250 2.7900 ;
        RECT  8.6650 2.1800 8.7850 2.7900 ;
        RECT  6.9350 1.8800 7.0550 2.7900 ;
        RECT  6.8150 1.8800 7.0550 2.0000 ;
        RECT  4.7750 1.7000 4.8950 2.7900 ;
        RECT  4.6550 1.7000 4.8950 1.9300 ;
        RECT  2.7150 1.9200 2.8350 2.7900 ;
        RECT  1.8150 1.4700 1.9350 2.7900 ;
        RECT  0.9750 1.3400 1.0950 2.7900 ;
        RECT  0.1350 1.3400 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.3850 0.8200 13.3650 0.8200 13.3650 1.6800 13.2850 1.6800 13.2850 1.8000
                 13.1650 1.8000 13.1650 1.6650 12.1850 1.6650 12.1850 1.2400 12.3050 1.2400
                 12.3050 1.5450 13.2450 1.5450 13.2450 0.7000 13.2650 0.7000 13.2650 0.5800
                 13.3850 0.5800 ;
        POLYGON  12.3250 0.8500 11.6050 0.8500 11.6050 1.5300 12.0650 1.5300 12.0650 2.2100
                 11.9450 2.2100 11.9450 1.6500 10.2650 1.6500 10.2650 1.6800 9.9650 1.6800
                 9.9650 2.0100 9.8450 2.0100 9.8450 1.5600 10.1450 1.5600 10.1450 0.8200 10.0050 0.8200
                 10.0050 0.7000 10.2650 0.7000 10.2650 1.5300 11.4850 1.5300 11.4850 0.7300
                 12.2050 0.7300 12.2050 0.5900 12.3250 0.5900 ;
        POLYGON  11.3650 1.0900 11.1250 1.0900 11.1250 0.8800 11.0050 0.8800 11.0050 0.5300
                 10.7400 0.5300 10.7400 0.5200 9.2700 0.5200 9.2700 0.8400 9.0050 0.8400 9.0050 0.8700
                 8.2850 0.8700 8.2850 0.5200 7.6100 0.5200 7.6100 0.8000 7.7750 0.8000 7.7750 1.5800
                 7.6550 1.5800 7.6550 0.9200 7.4900 0.9200 7.4900 0.4000 8.4050 0.4000 8.4050 0.7500
                 8.8850 0.7500 8.8850 0.7200 9.1500 0.7200 9.1500 0.4000 10.8600 0.4000 10.8600 0.4100
                 11.1250 0.4100 11.1250 0.7600 11.2450 0.7600 11.2450 0.9700 11.3650 0.9700 ;
        POLYGON  10.9450 2.2500 9.6050 2.2500 9.6050 1.4400 9.3650 1.4400 9.3650 1.2000 9.4850 1.2000
                 9.4850 1.3200 9.9050 1.3200 9.9050 0.9800 10.0250 0.9800 10.0250 1.4400 9.7250 1.4400
                 9.7250 2.1300 10.8250 2.1300 10.8250 1.7700 10.9450 1.7700 ;
        POLYGON  10.8650 0.7700 10.6250 0.7700 10.6250 1.0900 10.3850 1.0900 10.3850 0.9700
                 10.5050 0.9700 10.5050 0.6500 10.8650 0.6500 ;
        POLYGON  9.7650 1.0800 9.2450 1.0800 9.2450 1.5600 9.4850 1.5600 9.4850 2.2100 9.3650 2.2100
                 9.3650 1.6800 9.2450 1.6800 9.2450 2.0600 7.1750 2.0600 7.1750 1.7600 6.1150 1.7600
                 6.1150 1.9900 5.9950 1.9900 5.9950 1.4700 6.0950 1.4700 6.0950 0.7200 5.9950 0.7200
                 5.9950 0.6000 6.2350 0.6000 6.2350 0.7200 6.2150 0.7200 6.2150 1.6400 7.2950 1.6400
                 7.2950 1.9400 9.1250 1.9400 9.1250 0.9600 9.6450 0.9600 9.6450 0.6400 9.7650 0.6400 ;
        POLYGON  8.3050 1.8200 7.4150 1.8200 7.4150 1.5200 6.6950 1.5200 6.6950 1.2800 6.6550 1.2800
                 6.6550 1.0000 6.7750 1.0000 6.7750 1.1600 6.8150 1.1600 6.8150 1.4000 7.5350 1.4000
                 7.5350 1.7000 7.8950 1.7000 7.8950 0.7900 8.0450 0.7900 8.0450 0.6400 8.1650 0.6400
                 8.1650 0.9100 8.0150 0.9100 8.0150 1.5600 8.3050 1.5600 ;
        POLYGON  6.7100 0.8100 6.5350 0.8100 6.5350 1.4000 6.5750 1.4000 6.5750 1.5200 6.3350 1.5200
                 6.3350 1.4000 6.4150 1.4000 6.4150 0.6900 6.5900 0.6900 6.5900 0.5700 6.3550 0.5700
                 6.3550 0.4800 5.8750 0.4800 5.8750 1.1100 5.9750 1.1100 5.9750 1.3500 5.8550 1.3500
                 5.8550 1.2300 5.7550 1.2300 5.7550 0.4800 5.2750 0.4800 5.2750 0.8600 5.3950 0.8600
                 5.3950 1.1000 5.1550 1.1000 5.1550 0.8500 4.4150 0.8500 4.4150 0.4800 3.9350 0.4800
                 3.9350 0.8600 3.9750 0.8600 3.9750 1.1000 3.8150 1.1000 3.8150 0.4800 3.3350 0.4800
                 3.3350 0.8400 3.3950 0.8400 3.3950 1.3200 3.2750 1.3200 3.2750 0.9600 3.2150 0.9600
                 3.2150 0.3600 4.5350 0.3600 4.5350 0.7300 5.1550 0.7300 5.1550 0.3600 6.4750 0.3600
                 6.4750 0.4500 6.7100 0.4500 ;
        POLYGON  6.6950 2.2300 5.1300 2.2300 5.1300 1.5800 4.5350 1.5800 4.5350 2.2300 3.2650 2.2300
                 3.2650 1.8000 2.7350 1.8000 2.7350 1.3900 2.3550 1.3900 2.3550 1.9900 2.2350 1.9900
                 2.2350 1.5100 2.1550 1.5100 2.1550 1.2000 1.6350 1.2000 1.6350 1.0800 2.1550 1.0800
                 2.1550 0.6700 2.2350 0.6700 2.2350 0.5400 2.3550 0.5400 2.3550 0.7900 2.2750 0.7900
                 2.2750 1.2700 2.7350 1.2700 2.7350 1.1500 2.8550 1.1500 2.8550 1.6800 3.3850 1.6800
                 3.3850 2.1100 4.4150 2.1100 4.4150 1.4600 5.2500 1.4600 5.2500 2.1100 6.6950 2.1100 ;
        POLYGON  5.6350 1.9900 5.5150 1.9900 5.5150 1.3400 4.5750 1.3400 4.5750 1.3300 4.4550 1.3300
                 4.4550 1.2100 4.6950 1.2100 4.6950 1.2200 5.5150 1.2200 5.5150 0.7200 5.3950 0.7200
                 5.3950 0.6000 5.6350 0.6000 ;
        POLYGON  5.0350 1.0900 4.2950 1.0900 4.2950 1.9900 4.1750 1.9900 4.1750 0.7200 4.0550 0.7200
                 4.0550 0.6000 4.2950 0.6000 4.2950 0.9700 5.0350 0.9700 ;
        POLYGON  3.6950 0.7200 3.6350 0.7200 3.6350 1.9900 3.5150 1.9900 3.5150 1.5600 2.9750 1.5600
                 2.9750 1.0300 2.5150 1.0300 2.5150 1.1500 2.3950 1.1500 2.3950 0.9100 3.0950 0.9100
                 3.0950 1.4400 3.5150 1.4400 3.5150 0.7200 3.4550 0.7200 3.4550 0.6000 3.6950 0.6000 ;
    END
END SEDFFHQX4

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3700 0.7600 1.4900 1.1500 ;
        RECT  0.6300 0.7600 1.4900 0.8800 ;
        RECT  0.3050 1.2300 0.7500 1.3500 ;
        RECT  0.6300 0.7600 0.7500 1.3500 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.0300 1.0900 1.5000 ;
        RECT  0.9500 1.0000 1.0700 1.5000 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9400 2.8850 1.2100 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4600 1.0300 4.5800 1.4800 ;
        RECT  4.4200 1.0300 4.5800 1.4600 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0800 1.0800 11.2750 1.4350 ;
        RECT  11.0800 1.0750 11.2400 1.4350 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0300 1.5800 5.3400 1.7000 ;
        RECT  5.0000 0.6800 5.2400 0.8000 ;
        RECT  5.0300 0.6800 5.1500 1.7000 ;
        RECT  5.0000 0.6800 5.1500 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  10.7600 -0.1800 10.8800 0.7150 ;
        RECT  8.7700 -0.1800 9.0100 0.3900 ;
        RECT  6.9700 0.4600 7.2100 0.5800 ;
        RECT  6.9700 -0.1800 7.0900 0.5800 ;
        RECT  5.4800 -0.1800 5.7200 0.3200 ;
        RECT  4.5200 -0.1800 4.6400 0.6700 ;
        RECT  2.3500 0.4600 2.5900 0.5800 ;
        RECT  2.3500 -0.1800 2.4700 0.5800 ;
        RECT  0.8700 -0.1800 0.9900 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  10.8000 1.7950 10.9200 2.7900 ;
        RECT  8.5700 2.2500 8.8100 2.7900 ;
        RECT  6.8500 1.4700 6.9700 2.7900 ;
        RECT  5.5800 2.0600 5.8200 2.1800 ;
        RECT  5.5800 2.0600 5.7000 2.7900 ;
        RECT  4.7400 2.0600 4.8600 2.7900 ;
        RECT  4.6200 2.0600 4.8600 2.1800 ;
        RECT  2.4100 1.5700 2.5300 2.7900 ;
        RECT  0.8100 1.8600 0.9300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.4000 1.8550 11.1600 1.8550 11.1600 1.6750 10.6800 1.6750 10.6800 2.2500
                 9.1300 2.2500 9.1300 2.1300 8.1900 2.1300 8.1900 2.2500 7.8300 2.2500 7.8300 2.1300
                 8.0700 2.1300 8.0700 2.0100 9.3550 2.0100 9.3550 2.1300 10.5600 2.1300 10.5600 1.5550
                 10.8400 1.5550 10.8400 0.9550 10.7200 0.9550 10.7200 1.0750 10.6000 1.0750
                 10.6000 0.8350 11.1800 0.8350 11.1800 0.4750 11.3000 0.4750 11.3000 0.9550
                 10.9600 0.9550 10.9600 1.5550 11.2800 1.5550 11.2800 1.7350 11.4000 1.7350 ;
        POLYGON  10.4600 0.7150 10.4400 0.7150 10.4400 2.0100 9.6300 2.0100 9.6300 1.8900 7.8500 1.8900
                 7.8500 1.3300 7.4500 1.3300 7.4500 1.2100 7.8500 1.2100 7.8500 0.9900 8.2700 0.9900
                 8.2700 1.1100 7.9700 1.1100 7.9700 1.7700 9.6300 1.7700 9.6300 1.3300 9.5300 1.3300
                 9.5300 1.2100 9.7700 1.2100 9.7700 1.3300 9.7500 1.3300 9.7500 1.8900 10.3200 1.8900
                 10.3200 0.5950 10.3400 0.5950 10.3400 0.4750 10.4600 0.4750 ;
        POLYGON  10.1100 1.7700 9.8700 1.7700 9.8700 1.5300 9.9500 1.5300 9.9500 0.4800 9.2500 0.4800
                 9.2500 0.6300 8.5300 0.6300 8.5300 0.4800 7.4900 0.4800 7.4900 0.8200 6.7300 0.8200
                 6.7300 0.5300 6.0550 0.5300 6.0550 0.5600 4.8800 0.5600 4.8800 0.9100 4.1450 0.9100
                 4.1450 0.8600 4.0000 0.8600 4.0000 1.7700 3.8800 1.7700 3.8800 0.6200 4.0000 0.6200
                 4.0000 0.7400 4.2650 0.7400 4.2650 0.7900 4.7600 0.7900 4.7600 0.4400 5.9350 0.4400
                 5.9350 0.4100 6.8500 0.4100 6.8500 0.7000 7.3700 0.7000 7.3700 0.3600 8.6500 0.3600
                 8.6500 0.5100 9.1300 0.5100 9.1300 0.3600 10.0700 0.3600 10.0700 1.5300 10.1100 1.5300 ;
        POLYGON  9.7100 0.7200 9.5900 0.7200 9.5900 1.0900 9.4100 1.0900 9.4100 1.5300 9.5100 1.5300
                 9.5100 1.6500 9.2700 1.6500 9.2700 1.5300 9.2900 1.5300 9.2900 1.3600 8.6300 1.3600
                 8.6300 1.1200 8.7500 1.1200 8.7500 1.2400 9.2900 1.2400 9.2900 0.9700 9.4700 0.9700
                 9.4700 0.6000 9.7100 0.6000 ;
        POLYGON  9.0700 1.1200 8.9500 1.1200 8.9500 1.0000 8.5100 1.0000 8.5100 1.6500 8.0900 1.6500
                 8.0900 1.5300 8.3900 1.5300 8.3900 0.8700 8.1700 0.8700 8.1700 0.6000 8.4100 0.6000
                 8.4100 0.7500 8.5100 0.7500 8.5100 0.8800 9.0700 0.8800 ;
        POLYGON  7.9900 0.7200 7.7300 0.7200 7.7300 1.0600 7.3300 1.0600 7.3300 1.4500 7.7300 1.4500
                 7.7300 1.9900 7.6100 1.9900 7.6100 1.5700 7.2100 1.5700 7.2100 1.3500 6.6100 1.3500
                 6.6100 1.3300 6.4900 1.3300 6.4900 1.2100 6.7300 1.2100 6.7300 1.2300 7.2100 1.2300
                 7.2100 0.9400 7.6100 0.9400 7.6100 0.6000 7.9900 0.6000 ;
        POLYGON  7.0900 1.1100 6.8500 1.1100 6.8500 1.0900 6.3700 1.0900 6.3700 1.4700 6.5500 1.4700
                 6.5500 1.7800 6.4300 1.7800 6.4300 1.5900 6.2500 1.5900 6.2500 1.2100 6.1800 1.2100
                 6.1800 0.9700 6.2500 0.9700 6.2500 0.9200 6.3700 0.9200 6.3700 0.6500 6.6100 0.6500
                 6.6100 0.9700 6.9700 0.9700 6.9700 0.9900 7.0900 0.9900 ;
        POLYGON  6.2400 2.1700 6.1200 2.1700 6.1200 2.0500 5.9400 2.0500 5.9400 1.9400 4.4800 1.9400
                 4.4800 2.2500 2.6500 2.2500 2.6500 1.4500 2.2700 1.4500 2.2700 1.2100 2.3900 1.2100
                 2.3900 1.3300 2.7700 1.3300 2.7700 2.1300 4.3600 2.1300 4.3600 1.8200 5.9400 1.8200
                 5.9400 0.6800 6.2000 0.6800 6.2000 0.8000 6.0600 0.8000 6.0600 1.8200 6.2400 1.8200 ;
        POLYGON  4.2400 2.0100 2.8900 2.0100 2.8900 1.3300 3.0050 1.3300 3.0050 0.7700 2.9500 0.7700
                 2.9500 0.6500 3.1900 0.6500 3.1900 0.7700 3.1250 0.7700 3.1250 1.4500 3.0100 1.4500
                 3.0100 1.8900 3.6400 1.8900 3.6400 1.2000 3.5600 1.2000 3.5600 0.9600 3.7600 0.9600
                 3.7600 1.8900 4.1200 1.8900 4.1200 1.2000 4.2400 1.2000 ;
        POLYGON  3.5200 0.7700 3.4400 0.7700 3.4400 1.5200 3.5200 1.5200 3.5200 1.7700 3.4000 1.7700
                 3.4000 1.6400 3.3200 1.6400 3.3200 0.6500 3.4000 0.6500 3.4000 0.5300 2.8300 0.5300
                 2.8300 0.8200 1.7700 0.8200 1.7700 0.8300 1.7300 0.8300 1.7300 1.6600 1.5700 1.6600
                 1.5700 2.0100 1.4500 2.0100 1.4500 1.5400 1.6100 1.5400 1.6100 0.7100 1.6500 0.7100
                 1.6500 0.5900 1.7700 0.5900 1.7700 0.7000 2.7100 0.7000 2.7100 0.4100 3.5200 0.4100 ;
        POLYGON  2.0900 1.0900 1.9700 1.0900 1.9700 2.2500 1.2100 2.2500 1.2100 1.7400 0.4500 1.7400
                 0.4500 1.8600 0.3300 1.8600 0.3300 1.7400 0.0650 1.7400 0.0650 0.9900 0.3900 0.9900
                 0.3900 0.5900 0.5100 0.5900 0.5100 1.1100 0.1850 1.1100 0.1850 1.6200 1.2100 1.6200
                 1.2100 1.3000 1.4900 1.3000 1.4900 1.4200 1.3300 1.4200 1.3300 2.1300 1.8500 2.1300
                 1.8500 0.9700 2.0900 0.9700 ;
    END
END SEDFFHQX2

MACRO SEDFFHQX1
    CLASS CORE ;
    FOREIGN SEDFFHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3300 0.7600 1.4500 1.1500 ;
        RECT  0.5900 0.7600 1.4500 0.8800 ;
        RECT  0.4450 1.0700 0.7100 1.1900 ;
        RECT  0.5900 0.7600 0.7100 1.1900 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        RECT  0.4450 1.0700 0.5650 1.3800 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9100 1.0200 1.0900 1.4400 ;
        RECT  0.9100 1.0000 1.0300 1.4400 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9400 2.8850 1.1650 ;
        RECT  2.7100 0.9400 2.8300 1.3400 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3650 1.2250 4.6250 1.4600 ;
        RECT  4.3200 1.1300 4.5600 1.3450 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.8000 1.0300 10.9500 1.5000 ;
        RECT  10.8000 1.0300 10.9200 1.5300 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9000 0.6800 6.0200 1.0250 ;
        RECT  5.8950 0.9050 6.0150 1.9900 ;
        RECT  5.5800 1.0250 6.0150 1.1450 ;
        RECT  5.5800 0.8850 5.7300 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.6150 -0.1800 10.7350 0.6700 ;
        RECT  8.6250 0.4300 8.8650 0.5500 ;
        RECT  8.6250 -0.1800 8.7450 0.5500 ;
        RECT  6.9050 0.4100 7.1450 0.5300 ;
        RECT  6.9050 -0.1800 7.0250 0.5300 ;
        RECT  5.3600 -0.1800 5.6000 0.3200 ;
        RECT  4.4600 -0.1800 4.5800 0.6400 ;
        RECT  2.3100 0.4600 2.5500 0.5800 ;
        RECT  2.3100 -0.1800 2.4300 0.5800 ;
        RECT  0.8300 -0.1800 0.9500 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.6350 1.8900 10.7550 2.7900 ;
        RECT  8.4050 2.2500 8.6450 2.7900 ;
        RECT  6.8050 1.4900 6.9250 2.7900 ;
        RECT  5.4750 1.3400 5.5950 2.7900 ;
        RECT  4.5400 1.9000 4.6600 2.7900 ;
        RECT  2.2100 1.7000 2.3300 2.7900 ;
        RECT  0.7700 1.8000 0.8900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.2350 1.9500 10.9950 1.9500 10.9950 1.7700 10.5150 1.7700 10.5150 2.2500
                 8.9650 2.2500 8.9650 2.1300 8.0250 2.1300 8.0250 2.2500 7.6650 2.2500 7.6650 2.1300
                 7.9050 2.1300 7.9050 2.0100 9.0850 2.0100 9.0850 2.1300 10.3950 2.1300 10.3950 1.6500
                 10.5600 1.6500 10.5600 1.0300 10.4550 1.0300 10.4550 0.7900 10.8550 0.7900
                 10.8550 0.6700 11.0350 0.6700 11.0350 0.4300 11.1550 0.4300 11.1550 0.7900
                 10.9750 0.7900 10.9750 0.9100 10.6800 0.9100 10.6800 1.6500 11.1150 1.6500
                 11.1150 1.8300 11.2350 1.8300 ;
        POLYGON  10.3150 0.6700 10.2750 0.6700 10.2750 2.0100 9.4650 2.0100 9.4650 1.8900 7.6850 1.8900
                 7.6850 1.2500 7.4650 1.2500 7.4650 1.3700 7.3450 1.3700 7.3450 1.1300 7.9050 1.1300
                 7.9050 0.8600 8.0250 0.8600 8.0250 1.2500 7.8050 1.2500 7.8050 1.7700 9.4650 1.7700
                 9.4650 1.3300 9.3450 1.3300 9.3450 1.2100 9.5850 1.2100 9.5850 1.8900 10.1550 1.8900
                 10.1550 0.5500 10.1950 0.5500 10.1950 0.4300 10.3150 0.4300 ;
        POLYGON  9.9450 1.7700 9.7050 1.7700 9.7050 1.5300 9.8050 1.5300 9.8050 0.4800 9.1300 0.4800
                 9.1300 0.7900 8.3850 0.7900 8.3850 0.4800 7.3850 0.4800 7.3850 0.7700 6.6650 0.7700
                 6.6650 0.4800 6.1450 0.4800 6.1450 0.5600 4.8200 0.5600 4.8200 0.8800 4.0850 0.8800
                 4.0850 0.8300 3.9400 0.8300 3.9400 1.7700 3.8200 1.7700 3.8200 0.5900 3.9400 0.5900
                 3.9400 0.7100 4.2050 0.7100 4.2050 0.7600 4.7000 0.7600 4.7000 0.4400 6.0250 0.4400
                 6.0250 0.3600 6.7850 0.3600 6.7850 0.6500 7.2650 0.6500 7.2650 0.3600 8.5050 0.3600
                 8.5050 0.6700 9.0100 0.6700 9.0100 0.3600 9.9250 0.3600 9.9250 1.5300 9.9450 1.5300 ;
        POLYGON  9.5650 0.7200 9.4450 0.7200 9.4450 1.0900 9.2250 1.0900 9.2250 1.5300 9.3450 1.5300
                 9.3450 1.6500 9.1050 1.6500 9.1050 1.3900 8.3850 1.3900 8.3850 1.1500 8.5050 1.1500
                 8.5050 1.2700 9.1050 1.2700 9.1050 0.9700 9.3250 0.9700 9.3250 0.6000 9.5650 0.6000 ;
        POLYGON  8.8450 1.1500 8.7250 1.1500 8.7250 1.0300 8.2650 1.0300 8.2650 1.6500 7.9250 1.6500
                 7.9250 1.5300 8.1450 1.5300 8.1450 0.7200 8.0250 0.7200 8.0250 0.6000 8.2650 0.6000
                 8.2650 0.9100 8.8450 0.9100 ;
        POLYGON  7.8450 0.7200 7.7250 0.7200 7.7250 1.0100 7.2250 1.0100 7.2250 1.4900 7.5650 1.4900
                 7.5650 1.9900 7.4450 1.9900 7.4450 1.6100 7.1050 1.6100 7.1050 1.3700 6.5250 1.3700
                 6.5250 1.1300 6.6450 1.1300 6.6450 1.2500 7.1050 1.2500 7.1050 0.8900 7.6050 0.8900
                 7.6050 0.6000 7.8450 0.6000 ;
        POLYGON  6.9850 1.1300 6.8650 1.1300 6.8650 1.0100 6.4050 1.0100 6.4050 1.9900 6.2850 1.9900
                 6.2850 1.2400 6.1400 1.2400 6.1400 0.8900 6.2850 0.8900 6.2850 0.6000 6.5450 0.6000
                 6.5450 0.7200 6.4050 0.7200 6.4050 0.8900 6.9850 0.8900 ;
        POLYGON  5.1750 1.7800 4.4200 1.7800 4.4200 2.2500 2.4500 2.2500 2.4500 1.5800 2.1900 1.5800
                 2.1900 1.2400 2.3100 1.2400 2.3100 1.4600 2.5700 1.4600 2.5700 2.1300 4.3000 2.1300
                 4.3000 1.6600 5.0550 1.6600 5.0550 1.2200 4.9400 1.2200 4.9400 0.6800 5.0600 0.6800
                 5.0600 1.1000 5.1750 1.1000 ;
        POLYGON  4.1800 2.0100 2.6900 2.0100 2.6900 1.4600 3.0050 1.4600 3.0050 0.7700 2.9100 0.7700
                 2.9100 0.6500 3.1500 0.6500 3.1500 0.7700 3.1250 0.7700 3.1250 1.5800 2.8100 1.5800
                 2.8100 1.8900 3.5800 1.8900 3.5800 1.1700 3.5200 1.1700 3.5200 0.9300 3.7000 0.9300
                 3.7000 1.8900 4.0600 1.8900 4.0600 1.1500 4.1800 1.1500 ;
        POLYGON  3.4800 0.7700 3.4000 0.7700 3.4000 1.4900 3.4600 1.4900 3.4600 1.7700 3.3400 1.7700
                 3.3400 1.6100 3.2800 1.6100 3.2800 0.6500 3.3600 0.6500 3.3600 0.5300 2.7900 0.5300
                 2.7900 0.8200 1.7300 0.8200 1.7300 0.8300 1.6900 0.8300 1.6900 2.0100 1.5700 2.0100
                 1.5700 0.7100 1.6100 0.7100 1.6100 0.5900 1.7300 0.5900 1.7300 0.7000 2.6700 0.7000
                 2.6700 0.4100 3.4800 0.4100 ;
        POLYGON  2.0500 1.0900 1.9300 1.0900 1.9300 2.2500 1.3300 2.2500 1.3300 1.8000 1.2100 1.8000
                 1.2100 1.6800 0.4100 1.6800 0.4100 1.8000 0.2900 1.8000 0.2900 1.6800 0.0650 1.6800
                 0.0650 0.8300 0.3500 0.8300 0.3500 0.5900 0.4700 0.5900 0.4700 0.9500 0.1850 0.9500
                 0.1850 1.5600 1.2100 1.5600 1.2100 1.3000 1.4500 1.3000 1.4500 1.4200 1.3300 1.4200
                 1.3300 1.6800 1.4500 1.6800 1.4500 2.1300 1.8100 2.1300 1.8100 0.9700 2.0500 0.9700 ;
    END
END SEDFFHQX1

MACRO SDFFXL
    CLASS CORE ;
    FOREIGN SDFFXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 1.4100 2.1500 1.5400 ;
        RECT  1.7550 1.5100 2.0150 1.6700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0300 1.0200 7.1500 1.2600 ;
        RECT  6.7400 1.0200 7.1500 1.1400 ;
        RECT  6.7400 0.8850 6.8900 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4250 1.2100 8.6850 1.4450 ;
        RECT  8.3050 1.2100 8.6850 1.4200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0500 0.9400 8.8100 1.0600 ;
        RECT  8.6900 0.8200 8.8100 1.0600 ;
        RECT  8.0500 0.9400 8.3950 1.0900 ;
        RECT  7.5100 1.2400 8.1700 1.3600 ;
        RECT  8.0500 0.8200 8.1700 1.3600 ;
        RECT  7.5100 1.2400 7.6300 1.4800 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4100 1.3200 1.5300 1.9100 ;
        RECT  1.3700 0.6800 1.4900 0.9600 ;
        RECT  1.3300 0.8400 1.4500 1.4400 ;
        RECT  1.2300 0.8850 1.4500 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        RECT  8.5300 -0.1800 8.6500 0.7000 ;
        RECT  7.2500 -0.1800 7.3700 0.7000 ;
        RECT  5.0800 0.4500 5.3200 0.5700 ;
        RECT  5.2000 -0.1800 5.3200 0.5700 ;
        RECT  3.2000 0.6700 3.4400 0.7900 ;
        RECT  3.2400 -0.1800 3.3600 0.7900 ;
        RECT  1.7900 -0.1800 1.9100 0.4000 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        RECT  8.5300 1.9200 8.6500 2.7900 ;
        RECT  7.0900 1.9200 7.2100 2.7900 ;
        RECT  5.0400 2.2300 5.1600 2.7900 ;
        RECT  3.3800 2.1700 3.6200 2.2900 ;
        RECT  3.3800 2.1700 3.5000 2.7900 ;
        RECT  1.8300 1.7900 1.9500 2.7900 ;
        RECT  0.5550 1.4600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.0700 2.0400 8.9500 2.0400 8.9500 1.6850 8.0900 1.6850 8.0900 1.6600 7.9700 1.6600
                 7.9700 1.5400 8.2100 1.5400 8.2100 1.5650 8.9500 1.5650 8.9500 0.4600 9.0700 0.4600 ;
        POLYGON  8.0100 0.7000 7.9300 0.7000 7.9300 1.1200 7.3900 1.1200 7.3900 1.6000 7.4500 1.6000
                 7.4500 1.7200 7.8500 1.7200 7.8500 2.0400 7.7300 2.0400 7.7300 1.8400 7.3300 1.8400
                 7.3300 1.7200 6.5400 1.7200 6.5400 1.8100 6.2200 1.8100 6.2200 1.6900 6.4200 1.6900
                 6.4200 0.8200 6.3800 0.8200 6.3800 0.7000 6.6200 0.7000 6.6200 0.8200 6.5400 0.8200
                 6.5400 1.6000 7.2700 1.6000 7.2700 1.0000 7.8100 1.0000 7.8100 0.5800 7.8900 0.5800
                 7.8900 0.4600 8.0100 0.4600 ;
        POLYGON  6.9500 0.7000 6.8300 0.7000 6.8300 0.5800 6.2600 0.5800 6.2600 1.0600 6.1000 1.0600
                 6.1000 1.3500 6.3000 1.3500 6.3000 1.4700 6.1000 1.4700 6.1000 1.9300 6.8500 1.9300
                 6.8500 2.0500 5.9800 2.0500 5.9800 0.9400 6.1400 0.9400 6.1400 0.5800 5.5600 0.5800
                 5.5600 0.8100 4.8400 0.8100 4.8400 0.5200 4.4800 0.5200 4.4800 1.1700 4.6000 1.1700
                 4.6000 1.2900 4.3600 1.2900 4.3600 0.4000 4.9600 0.4000 4.9600 0.6900 5.4400 0.6900
                 5.4400 0.4600 5.6200 0.4600 5.6200 0.3600 5.8600 0.3600 5.8600 0.4600 6.9500 0.4600 ;
        POLYGON  6.0200 0.8200 5.8600 0.8200 5.8600 1.8700 5.7400 1.8700 5.7400 1.4100 4.9600 1.4100
                 4.9600 1.2900 5.7400 1.2900 5.7400 0.7000 6.0200 0.7000 ;
        POLYGON  5.7800 2.2500 5.4300 2.2500 5.4300 2.1100 4.6000 2.1100 4.6000 2.2500 4.3600 2.2500
                 4.3600 2.1100 3.8400 2.1100 3.8400 2.0500 2.5150 2.0500 2.5150 2.0300 2.2500 2.0300
                 2.2500 1.6700 2.2700 1.6700 2.2700 0.7400 2.5100 0.7400 2.5100 0.8600 2.3900 0.8600
                 2.3900 1.7900 2.3700 1.7900 2.3700 1.9100 2.6350 1.9100 2.6350 1.9300 3.8400 1.9300
                 3.8400 1.2700 3.7600 1.2700 3.7600 1.1500 4.0000 1.1500 4.0000 1.2700 3.9600 1.2700
                 3.9600 1.9900 5.5500 1.9900 5.5500 2.1300 5.7800 2.1300 ;
        POLYGON  5.5200 1.1700 4.8400 1.1700 4.8400 1.7500 4.6800 1.7500 4.6800 1.8700 4.5600 1.8700
                 4.5600 1.6300 4.7200 1.6300 4.7200 1.0500 4.6000 1.0500 4.6000 0.6400 4.7200 0.6400
                 4.7200 0.9300 4.8400 0.9300 4.8400 1.0500 5.5200 1.0500 ;
        POLYGON  4.3200 1.8100 4.0800 1.8100 4.0800 1.6900 4.1200 1.6900 4.1200 0.8800 3.8750 0.8800
                 3.8750 1.0300 2.9600 1.0300 2.9600 0.4800 2.8800 0.4800 2.8800 0.3600 3.1200 0.3600
                 3.1200 0.4800 3.0800 0.4800 3.0800 0.9100 3.7550 0.9100 3.7550 0.7600 4.1200 0.7600
                 4.1200 0.6400 4.2400 0.6400 4.2400 1.6900 4.3200 1.6900 ;
        POLYGON  3.6400 1.3900 3.0200 1.3900 3.0200 1.6900 3.1400 1.6900 3.1400 1.8100 2.9000 1.8100
                 2.9000 1.2700 2.7200 1.2700 2.7200 0.7200 2.6300 0.7200 2.6300 0.6200 2.1500 0.6200
                 2.1500 1.2000 1.5700 1.2000 1.5700 1.0800 2.0300 1.0800 2.0300 0.5000 2.7500 0.5000
                 2.7500 0.6000 2.8400 0.6000 2.8400 1.1500 3.0200 1.1500 3.0200 1.2700 3.6400 1.2700 ;
        POLYGON  1.1000 0.9200 1.0950 0.9200 1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000
                 0.3750 1.0800 0.9750 1.0800 0.9750 0.8000 0.9800 0.8000 0.9800 0.6800 1.1000 0.6800 ;
    END
END SDFFXL

MACRO SDFFX4
    CLASS CORE ;
    FOREIGN SDFFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0900 1.2000 1.2100 1.4400 ;
        RECT  0.3600 1.2000 1.2100 1.3200 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        RECT  0.3900 1.0800 0.5100 1.4350 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7700 1.4400 0.8900 1.7600 ;
        RECT  0.6500 1.4650 0.8000 1.7900 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.9900 1.9600 1.4500 ;
        RECT  1.8400 0.9650 1.9600 1.4500 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.4550 2.5950 1.6700 ;
        RECT  2.2150 1.4550 2.5950 1.6450 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0250 0.7000 9.2250 0.8200 ;
        RECT  9.0850 1.4400 9.2050 2.2100 ;
        RECT  8.9050 1.4400 9.2050 1.5600 ;
        RECT  8.2200 1.3200 9.0250 1.4400 ;
        RECT  8.2450 0.7000 8.3650 2.2100 ;
        RECT  8.1900 1.1750 8.3650 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.9450 0.7000 11.1450 0.8200 ;
        RECT  10.7650 1.3200 10.8850 2.2100 ;
        RECT  9.9300 1.3200 10.8850 1.4400 ;
        RECT  9.9600 0.7000 10.0800 1.5600 ;
        RECT  9.9250 1.4400 10.0450 2.2100 ;
        RECT  9.9300 1.1750 10.0800 1.5600 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.5050 -0.1800 11.6250 0.6900 ;
        RECT  10.4250 -0.1800 10.6650 0.3400 ;
        RECT  9.4650 -0.1800 9.7050 0.3400 ;
        RECT  8.5050 -0.1800 8.7450 0.3400 ;
        RECT  7.5450 -0.1800 7.7850 0.3400 ;
        RECT  6.7050 -0.1800 6.8250 0.8600 ;
        RECT  4.9850 0.5500 5.2250 0.6700 ;
        RECT  4.9850 -0.1800 5.1050 0.6700 ;
        RECT  2.9350 -0.1800 3.0550 0.9200 ;
        RECT  1.9500 -0.1800 2.0700 0.8450 ;
        RECT  0.6150 -0.1800 0.7350 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.1850 1.5600 11.3050 2.7900 ;
        RECT  10.3450 1.5600 10.4650 2.7900 ;
        RECT  9.5050 1.5600 9.6250 2.7900 ;
        RECT  8.6650 1.5600 8.7850 2.7900 ;
        RECT  7.8250 1.5600 7.9450 2.7900 ;
        RECT  6.9250 1.5800 7.0450 2.7900 ;
        RECT  5.2250 1.7500 5.3450 2.7900 ;
        RECT  3.3300 2.2900 3.5700 2.7900 ;
        RECT  2.1300 2.0500 2.3700 2.1700 ;
        RECT  2.1300 2.0500 2.2500 2.7900 ;
        RECT  0.7100 1.9500 0.8300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.0450 0.8800 11.8650 0.8800 11.8650 1.4400 11.7250 1.4400 11.7250 2.2100
                 11.6050 2.2100 11.6050 1.4400 11.0050 1.4400 11.0050 1.3000 11.2450 1.3000
                 11.2450 1.3200 11.7450 1.3200 11.7450 0.7600 11.9250 0.7600 11.9250 0.6400
                 12.0450 0.6400 ;
        POLYGON  11.5850 1.2000 11.4650 1.2000 11.4650 0.9300 11.2650 0.9300 11.2650 0.5800
                 7.2450 0.5800 7.2450 0.7000 7.6050 0.7000 7.6050 1.2600 8.0700 1.2600 8.0700 1.3800
                 7.4650 1.3800 7.4650 2.1000 7.3450 2.1000 7.3450 1.3800 6.9650 1.3800 6.9650 1.4600
                 6.8450 1.4600 6.8450 1.2200 6.9650 1.2200 6.9650 1.2600 7.4850 1.2600 7.4850 0.8200
                 7.1250 0.8200 7.1250 0.4600 11.3850 0.4600 11.3850 0.8100 11.5850 0.8100 ;
        POLYGON  7.3650 1.1400 7.1250 1.1400 7.1250 1.1000 6.7250 1.1000 6.7250 1.7700 6.3850 1.7700
                 6.3850 1.8100 6.1450 1.8100 6.1450 1.6900 6.2650 1.6900 6.2650 1.6500 6.6050 1.6500
                 6.6050 1.1000 6.0650 1.1000 6.0650 0.6200 6.1850 0.6200 6.1850 0.9800 7.3650 0.9800 ;
        POLYGON  6.4850 1.5300 6.3650 1.5300 6.3650 1.3400 5.8250 1.3400 5.8250 0.5000 5.4650 0.5000
                 5.4650 0.9100 4.7450 0.9100 4.7450 0.5000 4.1050 0.5000 4.1050 1.2900 4.2250 1.2900
                 4.2250 1.4100 3.9850 1.4100 3.9850 0.5000 3.4750 0.5000 3.4750 0.8000 3.6250 0.8000
                 3.6250 1.7700 3.9550 1.7700 3.9550 1.8900 3.5050 1.8900 3.5050 0.9200 3.3550 0.9200
                 3.3550 0.3800 4.4250 0.3800 4.4250 0.3600 4.6650 0.3600 4.6650 0.3800 4.8650 0.3800
                 4.8650 0.7900 5.3450 0.7900 5.3450 0.3800 5.9450 0.3800 5.9450 1.2200 6.4850 1.2200 ;
        POLYGON  5.7650 1.8700 5.6450 1.8700 5.6450 1.7500 5.5850 1.7500 5.5850 1.4900 5.0250 1.4900
                 5.0250 1.3700 5.5850 1.3700 5.5850 0.6200 5.7050 0.6200 5.7050 1.6300 5.7650 1.6300 ;
        POLYGON  5.4650 1.1500 4.6250 1.1500 4.6250 1.6300 4.7050 1.6300 4.7050 1.8700 4.5850 1.8700
                 4.5850 1.7500 4.5050 1.7500 4.5050 0.8000 4.2850 0.8000 4.2850 0.6800 4.6250 0.6800
                 4.6250 1.0300 5.4650 1.0300 ;
        POLYGON  4.2850 2.1100 4.2700 2.1100 4.2700 2.1300 3.2100 2.1300 3.2100 2.2500 2.4900 2.2500
                 2.4900 1.9300 1.4700 1.9300 1.4700 2.0700 1.3500 2.0700 1.3500 1.9500 1.3300 1.9500
                 1.3300 0.8400 1.1900 0.8400 1.1900 0.7200 1.4500 0.7200 1.4500 1.8100 2.6100 1.8100
                 2.6100 2.1300 3.0900 2.1300 3.0900 2.0100 4.1500 2.0100 4.1500 1.9900 4.1650 1.9900
                 4.1650 1.6500 3.7450 1.6500 3.7450 0.6200 3.8650 0.6200 3.8650 1.5300 4.2850 1.5300 ;
        POLYGON  3.3850 1.2100 2.8500 1.2100 2.8500 1.8900 2.9700 1.8900 2.9700 2.0100 2.7300 2.0100
                 2.7300 1.1600 2.4300 1.1600 2.4300 0.6600 2.5500 0.6600 2.5500 1.0400 2.8500 1.0400
                 2.8500 1.0900 3.3850 1.0900 ;
        POLYGON  1.8100 1.6900 1.5700 1.6900 1.5700 0.6000 1.0050 0.6000 1.0050 0.6600 0.2550 0.6600
                 0.2550 0.9000 0.2400 0.9000 0.2400 1.5550 0.4100 1.5550 0.4100 2.0700 0.2900 2.0700
                 0.2900 1.6750 0.1200 1.6750 0.1200 0.7800 0.1350 0.7800 0.1350 0.5400 0.8850 0.5400
                 0.8850 0.4800 1.0300 0.4800 1.0300 0.3800 1.2700 0.3800 1.2700 0.4800 1.6900 0.4800
                 1.6900 1.5700 1.8100 1.5700 ;
    END
END SDFFX4

MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4050 1.2250 1.2850 1.3450 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        RECT  0.4050 1.2250 0.5250 1.4700 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.4650 1.0900 1.7850 ;
        RECT  0.6850 1.4650 1.0900 1.6150 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.5800 ;
        RECT  2.0050 1.2550 2.1250 1.6700 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0600 0.7400 7.1800 1.2600 ;
        RECT  7.0300 0.7400 7.1800 1.2000 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8300 1.1750 8.0500 1.4350 ;
        RECT  7.8300 0.7400 7.9500 2.0100 ;
        RECT  7.6500 0.7400 7.9500 0.8600 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.6100 0.7400 8.8500 0.8600 ;
        RECT  8.6700 0.7400 8.7900 2.0100 ;
        RECT  8.4800 0.8850 8.7900 1.1450 ;
        RECT  8.6100 0.7400 8.7900 1.1450 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.1500 -0.1800 9.2700 0.3800 ;
        RECT  8.1300 -0.1800 8.3700 0.3800 ;
        RECT  7.1700 -0.1800 7.4100 0.3800 ;
        RECT  5.8600 0.6800 6.1000 0.8000 ;
        RECT  5.8600 -0.1800 5.9800 0.8000 ;
        RECT  4.1400 -0.1800 4.3800 0.3200 ;
        RECT  1.9450 -0.1800 2.0650 0.8600 ;
        RECT  0.5450 0.6800 0.7850 0.8000 ;
        RECT  0.5450 -0.1800 0.6650 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  9.0900 1.3600 9.2100 2.7900 ;
        RECT  8.2500 1.3600 8.3700 2.7900 ;
        RECT  7.4100 1.3600 7.5300 2.7900 ;
        RECT  5.8950 2.1400 6.1350 2.2600 ;
        RECT  5.8950 2.1400 6.0150 2.7900 ;
        RECT  4.2550 2.2000 4.4950 2.7900 ;
        RECT  2.1450 2.1800 2.3850 2.3000 ;
        RECT  2.1450 2.1800 2.2650 2.7900 ;
        RECT  0.6650 1.9500 0.7850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.7850 0.8600 9.6650 0.8600 9.6650 1.1800 9.6300 1.1800 9.6300 1.6000 9.5100 1.6000
                 9.5100 1.1800 8.9100 1.1800 8.9100 1.0600 9.5450 1.0600 9.5450 0.7400 9.7850 0.7400 ;
        POLYGON  9.6500 0.5200 9.5300 0.5200 9.5300 0.6200 8.2900 0.6200 8.2900 1.2400 8.1700 1.2400
                 8.1700 0.6200 7.4950 0.6200 7.4950 1.0600 7.6150 1.0600 7.6150 1.1800 7.3750 1.1800
                 7.3750 0.6200 6.4600 0.6200 6.4600 0.7400 6.5350 0.7400 6.5350 1.6600 6.6150 1.6600
                 6.6150 1.7800 6.3750 1.7800 6.3750 1.6600 6.4150 1.6600 6.4150 1.4000 6.0150 1.4000
                 6.0150 1.5200 5.8950 1.5200 5.8950 1.2800 6.4150 1.2800 6.4150 0.8600 6.3400 0.8600
                 6.3400 0.5000 9.4100 0.5000 9.4100 0.4000 9.6500 0.4000 ;
        POLYGON  7.0500 2.0200 5.5250 2.0200 5.5250 2.0800 5.2950 2.0800 5.2950 2.2200 5.0550 2.2200
                 5.0550 2.0800 3.9350 2.0800 3.9350 2.2200 3.6950 2.2200 3.6950 2.1000 3.8150 2.1000
                 3.8150 1.9600 5.4050 1.9600 5.4050 1.9000 6.9300 1.9000 6.9300 1.5000 6.7900 1.5000
                 6.7900 0.8600 6.6700 0.8600 6.6700 0.7400 6.9100 0.7400 6.9100 1.3800 7.0500 1.3800 ;
        POLYGON  6.2950 1.1400 5.7750 1.1400 5.7750 1.7400 5.4350 1.7400 5.4350 1.7800 5.1950 1.7800
                 5.1950 1.6600 5.3150 1.6600 5.3150 1.6200 5.6550 1.6200 5.6550 1.1400 5.3400 1.1400
                 5.3400 0.8000 5.2200 0.8000 5.2200 0.6800 5.4600 0.6800 5.4600 1.0200 6.2950 1.0200 ;
        POLYGON  5.5350 1.5000 5.4150 1.5000 5.4150 1.3800 4.9800 1.3800 4.9800 1.2000 4.8750 1.2000
                 4.8750 0.9600 4.9800 0.9600 4.9800 0.5600 3.3200 0.5600 3.3200 1.2200 3.3800 1.2200
                 3.3800 1.3400 3.1400 1.3400 3.1400 1.2200 3.2000 1.2200 3.2000 0.5600 2.7200 0.5600
                 2.7200 0.6200 2.4850 0.6200 2.4850 0.7400 2.4900 0.7400 2.4900 1.7000 2.9850 1.7000
                 2.9850 2.0100 2.7450 2.0100 2.7450 1.8200 2.3700 1.8200 2.3700 0.8600 2.3650 0.8600
                 2.3650 0.5000 2.6000 0.5000 2.6000 0.4400 3.5800 0.4400 3.5800 0.3600 3.8200 0.3600
                 3.8200 0.4400 5.1000 0.4400 5.1000 1.2600 5.5350 1.2600 ;
        POLYGON  4.9150 1.8400 4.7950 1.8400 4.7950 1.6200 4.7400 1.6200 4.7400 1.4600 4.0550 1.4600
                 4.0550 1.3400 4.6350 1.3400 4.6350 0.8000 4.6200 0.8000 4.6200 0.6800 4.8600 0.6800
                 4.8600 0.8000 4.7550 0.8000 4.7550 1.3400 4.8600 1.3400 4.8600 1.5000 4.9150 1.5000 ;
        POLYGON  4.5150 1.1400 3.7350 1.1400 3.7350 1.8400 3.6150 1.8400 3.6150 0.8000 3.4400 0.8000
                 3.4400 0.6800 3.7350 0.6800 3.7350 1.0200 4.5150 1.0200 ;
        POLYGON  3.3150 2.2500 2.5050 2.2500 2.5050 2.0600 1.5250 2.0600 1.5250 2.0700 1.4050 2.0700
                 1.4050 0.8000 1.1850 0.8000 1.1850 0.6800 1.5250 0.6800 1.5250 1.9400 2.6250 1.9400
                 2.6250 2.1300 3.1950 2.1300 3.1950 1.5800 2.9000 1.5800 2.9000 0.8000 2.8400 0.8000
                 2.8400 0.6800 3.0800 0.6800 3.0800 0.8000 3.0200 0.8000 3.0200 1.4600 3.3150 1.4600 ;
        POLYGON  1.7650 1.7500 1.6450 1.7500 1.6450 0.5600 1.0250 0.5600 1.0250 1.0400 0.1850 1.0400
                 0.1850 1.5900 0.3650 1.5900 0.3650 2.0700 0.2450 2.0700 0.2450 1.7100 0.0650 1.7100
                 0.0650 0.7400 0.1850 0.7400 0.1850 0.6200 0.3050 0.6200 0.3050 0.9200 0.9050 0.9200
                 0.9050 0.4400 1.0450 0.4400 1.0450 0.3600 1.2850 0.3600 1.2850 0.4400 1.7650 0.4400 ;
    END
END SDFFX2

MACRO SDFFX1
    CLASS CORE ;
    FOREIGN SDFFX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1300 1.2200 2.2500 1.4600 ;
        RECT  1.7550 1.5200 2.1500 1.6700 ;
        RECT  2.0300 1.3400 2.1500 1.6700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9150 1.2900 7.0350 1.5300 ;
        RECT  6.7400 1.2900 7.0350 1.4350 ;
        RECT  6.7400 1.1750 6.8900 1.4350 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1150 1.2300 8.3950 1.4700 ;
        RECT  8.1350 1.2100 8.3950 1.4700 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4250 0.9400 8.6850 1.0900 ;
        RECT  8.4750 0.8500 8.5950 1.0900 ;
        RECT  7.5150 0.9500 8.6850 1.0700 ;
        RECT  7.7550 0.8700 7.9950 1.0700 ;
        RECT  7.3950 1.4100 7.6350 1.5300 ;
        RECT  7.5150 0.9500 7.6350 1.5300 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 0.8850 1.6700 1.1450 ;
        RECT  1.4550 0.8850 1.5750 2.2100 ;
        RECT  1.3950 0.6800 1.5150 1.0250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.3150 -0.1800 8.4350 0.7300 ;
        RECT  7.0350 -0.1800 7.1550 0.7300 ;
        RECT  4.8450 -0.1800 5.0850 0.3200 ;
        RECT  3.2250 -0.1800 3.4650 0.3200 ;
        RECT  1.7550 0.5500 1.9950 0.6700 ;
        RECT  1.7550 -0.1800 1.8750 0.6700 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.3150 1.8300 8.4350 2.7900 ;
        RECT  6.8350 1.8900 7.0750 2.0100 ;
        RECT  6.8350 1.8900 6.9550 2.7900 ;
        RECT  4.8650 2.1600 4.9850 2.7900 ;
        RECT  3.2050 2.1600 3.4450 2.2800 ;
        RECT  3.2050 2.1600 3.3250 2.7900 ;
        RECT  1.8750 1.7900 1.9950 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.9250 1.8300 8.8550 1.8300 8.8550 1.9500 8.7350 1.9500 8.7350 1.7100 7.8750 1.7100
                 7.8750 1.3100 7.7550 1.3100 7.7550 1.1900 7.9950 1.1900 7.9950 1.5900 8.8050 1.5900
                 8.8050 0.8200 8.7350 0.8200 8.7350 0.4900 8.8550 0.4900 8.8550 0.7000 8.9250 0.7000 ;
        POLYGON  7.7950 0.7500 7.3950 0.7500 7.3950 1.2900 7.2750 1.2900 7.2750 1.6500 7.6550 1.6500
                 7.6550 1.9500 7.5350 1.9500 7.5350 1.7700 6.1650 1.7700 6.1650 1.8800 6.0450 1.8800
                 6.0450 1.6400 6.1450 1.6400 6.1450 0.6600 6.2650 0.6600 6.2650 1.6500 7.1550 1.6500
                 7.1550 1.1700 7.2750 1.1700 7.2750 0.6300 7.6750 0.6300 7.6750 0.4900 7.7950 0.4900 ;
        POLYGON  6.7950 0.6700 6.5550 0.6700 6.5550 0.5400 6.0250 0.5400 6.0250 1.0800 5.9250 1.0800
                 5.9250 1.2800 6.0050 1.2800 6.0050 1.5200 5.9250 1.5200 5.9250 2.0000 6.3750 2.0000
                 6.3750 1.8900 6.6150 1.8900 6.6150 2.0100 6.4950 2.0100 6.4950 2.1200 5.8050 2.1200
                 5.8050 0.9600 5.9050 0.9600 5.9050 0.5400 5.3800 0.5400 5.3800 0.5600 4.3250 0.5600
                 4.3250 1.2200 4.2050 1.2200 4.2050 0.4400 5.2600 0.4400 5.2600 0.4200 5.4050 0.4200
                 5.4050 0.4000 5.6450 0.4000 5.6450 0.4200 6.6750 0.4200 6.6750 0.5500 6.7950 0.5500 ;
        POLYGON  5.7850 0.8400 5.6850 0.8400 5.6850 1.8600 5.5650 1.8600 5.5650 1.4800 4.7250 1.4800
                 4.7250 1.3600 5.5650 1.3600 5.5650 0.8400 5.5450 0.8400 5.5450 0.7200 5.7850 0.7200 ;
        POLYGON  5.6050 2.2400 5.3250 2.2400 5.3250 2.0400 4.5950 2.0400 4.5950 2.1000 4.4250 2.1000
                 4.4250 2.2400 4.1850 2.2400 4.1850 2.1000 3.6800 2.1000 3.6800 2.0400 2.3550 2.0400
                 2.3550 1.6800 2.3700 1.6800 2.3700 1.1000 2.3550 1.1000 2.3550 0.6800 2.4750 0.6800
                 2.4750 0.9800 2.4900 0.9800 2.4900 1.8000 2.4750 1.8000 2.4750 1.9200 3.6800 1.9200
                 3.6800 1.1600 3.6050 1.1600 3.6050 1.0400 3.8450 1.0400 3.8450 1.1600 3.8000 1.1600
                 3.8000 1.9800 4.4750 1.9800 4.4750 1.9200 5.4450 1.9200 5.4450 2.1200 5.6050 2.1200 ;
        POLYGON  5.1850 1.2200 4.5650 1.2200 4.5650 1.8000 4.3250 1.8000 4.3250 1.6800 4.4450 1.6800
                 4.4450 0.7200 4.6850 0.7200 4.6850 0.8400 4.5650 0.8400 4.5650 1.1000 5.0650 1.1000
                 5.0650 0.9800 5.1850 0.9800 ;
        POLYGON  4.0850 1.8600 3.9650 1.8600 3.9650 0.9000 3.9250 0.9000 3.9250 0.6600 2.9850 0.6600
                 2.9850 0.5000 2.8450 0.5000 2.8450 0.3800 3.1050 0.3800 3.1050 0.5400 4.0450 0.5400
                 4.0450 0.7800 4.0850 0.7800 ;
        POLYGON  3.4850 1.2400 2.8650 1.2400 2.8650 1.6800 2.9650 1.6800 2.9650 1.8000 2.7250 1.8000
                 2.7250 1.6800 2.7450 1.6800 2.7450 0.7800 2.6050 0.7800 2.6050 0.5600 2.2350 0.5600
                 2.2350 0.9100 1.9100 0.9100 1.9100 1.2400 1.7900 1.2400 1.7900 0.7900 2.1150 0.7900
                 2.1150 0.4400 2.7250 0.4400 2.7250 0.6600 2.8650 0.6600 2.8650 1.1200 3.4850 1.1200 ;
        POLYGON  1.1550 1.5800 1.0350 1.5800 1.0350 1.3200 1.0050 1.3200 1.0050 1.2000 0.3750 1.2000
                 0.3750 1.0800 1.0050 1.0800 1.0050 0.6800 1.1250 0.6800 1.1250 1.2000 1.1550 1.2000 ;
    END
END SDFFX1

MACRO SDFFTRXL
    CLASS CORE ;
    FOREIGN SDFFTRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 1.4100 2.1450 1.5400 ;
        RECT  1.7550 1.5100 2.0150 1.6700 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8700 1.1600 7.0150 1.4000 ;
        RECT  6.7400 1.1750 6.9150 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7350 0.9400 8.9750 1.3000 ;
        RECT  8.7150 0.9400 8.9750 1.0900 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.1550 0.9400 9.5550 1.1700 ;
        RECT  9.1550 0.9400 9.2750 1.3500 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6750 0.9600 10.1350 1.1500 ;
        RECT  9.8750 0.9350 10.1350 1.1500 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4050 1.3200 1.5250 1.9100 ;
        RECT  1.3650 0.6800 1.4850 0.9600 ;
        RECT  1.2300 1.1750 1.4450 1.4350 ;
        RECT  1.3250 0.8400 1.4450 1.4400 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  9.0150 -0.1800 9.1350 0.8200 ;
        RECT  6.9950 -0.1800 7.1150 0.8400 ;
        RECT  4.9450 -0.1800 5.1850 0.3400 ;
        RECT  3.2450 -0.1800 3.4850 0.3400 ;
        RECT  1.7850 -0.1800 1.9050 0.4000 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  9.8550 1.5800 9.9750 2.7900 ;
        RECT  8.9550 2.0600 9.0750 2.7900 ;
        RECT  6.8950 1.8400 7.0150 2.7900 ;
        RECT  4.9050 2.1600 5.0250 2.7900 ;
        RECT  3.2450 2.1000 3.4850 2.2200 ;
        RECT  3.2450 2.1000 3.3650 2.7900 ;
        RECT  1.8250 1.7900 1.9450 2.7900 ;
        RECT  0.5550 1.4600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.3750 1.4600 9.5550 1.4600 9.5550 1.8300 9.1350 1.8300 9.1350 1.9400 8.0750 1.9400
                 8.0750 1.9600 7.9550 1.9600 7.9550 1.4400 8.2350 1.4400 8.2350 0.8400 8.1150 0.8400
                 8.1150 0.6000 8.2350 0.6000 8.2350 0.7200 8.3550 0.7200 8.3550 1.5600 8.0750 1.5600
                 8.0750 1.8200 9.0150 1.8200 9.0150 1.7100 9.4350 1.7100 9.4350 1.3400 10.2550 1.3400
                 10.2550 0.7600 9.5950 0.7600 9.5950 0.6400 10.3750 0.6400 ;
        POLYGON  8.7150 0.8200 8.5950 0.8200 8.5950 1.7000 8.4750 1.7000 8.4750 0.7000 8.5950 0.7000
                 8.5950 0.5800 8.4050 0.5800 8.4050 0.4800 7.9950 0.4800 7.9950 0.9800 8.1150 0.9800
                 8.1150 1.1000 7.9950 1.1000 7.9950 1.3200 7.4950 1.3200 7.4950 1.4800 7.3750 1.4800
                 7.3750 1.2000 7.8750 1.2000 7.8750 0.3600 8.5250 0.3600 8.5250 0.4600 8.7150 0.4600 ;
        POLYGON  7.7550 1.0800 7.2550 1.0800 7.2550 1.6000 7.6550 1.6000 7.6550 1.9600 7.5350 1.9600
                 7.5350 1.7200 6.2050 1.7200 6.2050 1.8400 6.0850 1.8400 6.0850 1.6000 6.1850 1.6000
                 6.1850 0.6800 6.3050 0.6800 6.3050 1.6000 7.1350 1.6000 7.1350 0.9600 7.6350 0.9600
                 7.6350 0.6000 7.7550 0.6000 ;
        POLYGON  6.6950 0.8400 6.5750 0.8400 6.5750 0.6000 6.4750 0.6000 6.4750 0.5600 6.0650 0.5600
                 6.0650 1.1000 5.9650 1.1000 5.9650 1.2400 6.0650 1.2400 6.0650 1.4800 5.9650 1.4800
                 5.9650 1.9600 6.4150 1.9600 6.4150 1.9000 6.6550 1.9000 6.6550 2.0200 6.5350 2.0200
                 6.5350 2.0800 5.8450 2.0800 5.8450 0.9800 5.9450 0.9800 5.9450 0.5600 5.4250 0.5600
                 5.4250 0.5800 4.7050 0.5800 4.7050 0.5600 4.3450 0.5600 4.3450 1.2600 4.2250 1.2600
                 4.2250 0.4400 4.8250 0.4400 4.8250 0.4600 5.3050 0.4600 5.3050 0.4400 5.4250 0.4400
                 5.4250 0.4000 5.6650 0.4000 5.6650 0.4400 6.5950 0.4400 6.5950 0.4800 6.6950 0.4800 ;
        POLYGON  5.8250 0.8600 5.7250 0.8600 5.7250 1.8000 5.6050 1.8000 5.6050 1.4400 4.8250 1.4400
                 4.8250 1.4200 4.7050 1.4200 4.7050 1.3000 4.9450 1.3000 4.9450 1.3200 5.6050 1.3200
                 5.6050 0.8600 5.5850 0.8600 5.5850 0.7400 5.8250 0.7400 ;
        POLYGON  5.6450 2.1800 5.4050 2.1800 5.4050 2.0400 4.3250 2.0400 4.3250 2.1800 4.0850 2.1800
                 4.0850 2.0400 3.6250 2.0400 3.6250 1.9800 2.2450 1.9800 2.2450 1.6700 2.2650 1.6700
                 2.2650 0.7400 2.5050 0.7400 2.5050 0.8600 2.3850 0.8600 2.3850 1.8600 3.6250 1.8600
                 3.6250 1.0600 3.8650 1.0600 3.8650 1.1800 3.7450 1.1800 3.7450 1.9200 5.5250 1.9200
                 5.5250 2.0600 5.6450 2.0600 ;
        POLYGON  5.3050 1.2000 5.0650 1.2000 5.0650 1.1800 4.5850 1.1800 4.5850 1.5000 4.5450 1.5000
                 4.5450 1.8000 4.4250 1.8000 4.4250 1.3800 4.4650 1.3800 4.4650 0.6800 4.5850 0.6800
                 4.5850 1.0600 5.1850 1.0600 5.1850 1.0800 5.3050 1.0800 ;
        POLYGON  4.1250 1.8000 4.0050 1.8000 4.0050 1.5000 3.9850 1.5000 3.9850 0.9200 3.9650 0.9200
                 3.9650 0.6800 3.0050 0.6800 3.0050 0.5200 2.8650 0.5200 2.8650 0.4000 3.1250 0.4000
                 3.1250 0.5600 4.0850 0.5600 4.0850 0.8000 4.1050 0.8000 4.1050 1.3800 4.1250 1.3800 ;
        POLYGON  3.5050 1.2600 2.8850 1.2600 2.8850 1.6200 3.0050 1.6200 3.0050 1.7400 2.7650 1.7400
                 2.7650 0.8000 2.6250 0.8000 2.6250 0.6200 2.1450 0.6200 2.1450 1.2000 1.5650 1.2000
                 1.5650 1.0800 2.0250 1.0800 2.0250 0.5000 2.7450 0.5000 2.7450 0.6800 2.8850 0.6800
                 2.8850 1.1400 3.5050 1.1400 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END SDFFTRXL

MACRO SDFFTRX4
    CLASS CORE ;
    FOREIGN SDFFTRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.3400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4050 1.1000 0.5250 1.3400 ;
        RECT  0.0700 1.1750 0.5250 1.2950 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0900 1.0400 1.2100 1.4300 ;
        RECT  0.8850 1.1900 1.2100 1.4100 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.2000 1.7250 1.4100 ;
        RECT  1.6050 1.0400 1.7250 1.4100 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.1750 3.4100 1.4350 ;
        RECT  3.1200 1.1750 3.4100 1.2950 ;
        RECT  3.1200 1.0550 3.2400 1.2950 ;
        END
    END SI
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 1.1750 3.7000 1.5350 ;
        RECT  3.5300 1.0000 3.6500 1.3650 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.1850 0.7200 10.3850 0.8400 ;
        RECT  10.2450 1.4400 10.3650 2.2100 ;
        RECT  10.0650 1.4400 10.3650 1.5600 ;
        RECT  9.3800 1.3200 10.1850 1.4400 ;
        RECT  9.4050 0.7200 9.5250 2.2100 ;
        RECT  9.3500 1.1750 9.5250 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.1050 0.7200 12.3050 0.8400 ;
        RECT  11.9250 1.3200 12.0450 2.2100 ;
        RECT  11.0900 1.3200 12.0450 1.4400 ;
        RECT  11.1200 0.7200 11.2400 1.5600 ;
        RECT  11.0850 1.4400 11.2050 2.2100 ;
        RECT  11.0900 1.1750 11.2400 1.5600 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.3400 0.1800 ;
        RECT  12.6650 -0.1800 12.7850 0.7100 ;
        RECT  11.5850 -0.1800 11.8250 0.3600 ;
        RECT  10.6250 -0.1800 10.8650 0.3600 ;
        RECT  9.6650 -0.1800 9.9050 0.3600 ;
        RECT  8.7050 -0.1800 8.9450 0.3600 ;
        RECT  7.8650 -0.1800 7.9850 0.9000 ;
        RECT  6.1450 -0.1800 6.3850 0.3200 ;
        RECT  4.2150 -0.1800 4.3350 0.9200 ;
        RECT  3.2200 -0.1800 3.3400 0.8800 ;
        RECT  1.2300 -0.1800 1.3500 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.3400 2.7900 ;
        RECT  12.3450 1.5800 12.4650 2.7900 ;
        RECT  11.5050 1.5600 11.6250 2.7900 ;
        RECT  10.6650 1.5600 10.7850 2.7900 ;
        RECT  9.8250 1.5600 9.9450 2.7900 ;
        RECT  8.9850 1.5600 9.1050 2.7900 ;
        RECT  8.0850 1.6200 8.2050 2.7900 ;
        RECT  6.2050 1.7400 6.3250 2.7900 ;
        RECT  4.3000 1.9800 4.4200 2.7900 ;
        RECT  3.2200 1.9400 3.3400 2.7900 ;
        RECT  1.2900 2.0100 1.4100 2.7900 ;
        RECT  0.3900 1.5900 0.5100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.2050 0.9000 13.0250 0.9000 13.0250 1.4600 12.8850 1.4600 12.8850 2.2100
                 12.7650 2.2100 12.7650 1.4600 12.1650 1.4600 12.1650 1.3000 12.4050 1.3000
                 12.4050 1.3400 12.9050 1.3400 12.9050 0.7800 13.0850 0.7800 13.0850 0.6600
                 13.2050 0.6600 ;
        POLYGON  12.7450 1.2200 12.6250 1.2200 12.6250 0.9500 12.4250 0.9500 12.4250 0.6000
                 8.9350 0.6000 8.9350 0.6600 8.4050 0.6600 8.4050 0.7800 8.7650 0.7800 8.7650 1.2800
                 9.2300 1.2800 9.2300 1.4000 8.6250 1.4000 8.6250 2.1400 8.5050 2.1400 8.5050 1.4000
                 8.1250 1.4000 8.1250 1.5000 8.0050 1.5000 8.0050 1.2600 8.1250 1.2600 8.1250 1.2800
                 8.6450 1.2800 8.6450 0.9000 8.2850 0.9000 8.2850 0.5400 8.8150 0.5400 8.8150 0.4800
                 12.5450 0.4800 12.5450 0.8300 12.7450 0.8300 ;
        POLYGON  8.5250 1.1600 8.2850 1.1600 8.2850 1.1400 7.8850 1.1400 7.8850 1.7600 7.5450 1.7600
                 7.5450 1.8000 7.3050 1.8000 7.3050 1.6800 7.4250 1.6800 7.4250 1.6400 7.7650 1.6400
                 7.7650 1.1400 7.2250 1.1400 7.2250 0.6600 7.3450 0.6600 7.3450 1.0200 8.5250 1.0200 ;
        POLYGON  7.6450 1.5200 7.5250 1.5200 7.5250 1.3800 6.9850 1.3800 6.9850 0.5400 6.6250 0.5400
                 6.6250 0.5600 5.9050 0.5600 5.9050 0.5400 5.3850 0.5400 5.3850 1.3600 5.4450 1.3600
                 5.4450 1.4800 5.2050 1.4800 5.2050 1.3600 5.2650 1.3600 5.2650 0.5400 4.8550 0.5400
                 4.8550 0.6800 4.7550 0.6800 4.7550 0.8000 4.8450 0.8000 4.8450 1.5800 4.7250 1.5800
                 4.7250 0.9200 4.6350 0.9200 4.6350 0.5600 4.7350 0.5600 4.7350 0.4200 5.6650 0.4200
                 5.6650 0.3800 5.9050 0.3800 5.9050 0.4200 6.0250 0.4200 6.0250 0.4400 6.5050 0.4400
                 6.5050 0.4200 7.1050 0.4200 7.1050 1.2600 7.6450 1.2600 ;
        POLYGON  6.8650 1.8600 6.7450 1.8600 6.7450 1.4800 6.0050 1.4800 6.0050 1.3600 6.7450 1.3600
                 6.7450 0.6600 6.8650 0.6600 ;
        POLYGON  6.6250 1.2400 5.6850 1.2400 5.6850 1.8600 5.5650 1.8600 5.5650 0.8400 5.5050 0.8400
                 5.5050 0.7200 5.7450 0.7200 5.7450 0.8400 5.6850 0.8400 5.6850 1.1200 6.6250 1.1200 ;
        POLYGON  5.2450 1.8600 4.1800 1.8600 4.1800 2.2400 3.4600 2.2400 3.4600 1.8200 2.9650 1.8200
                 2.9650 1.9400 2.7000 1.9400 2.7000 2.0600 2.5800 2.0600 2.5800 1.9400 2.4400 1.9400
                 2.4400 0.7000 2.7600 0.7000 2.7600 0.8200 2.5600 0.8200 2.5600 1.8200 2.8450 1.8200
                 2.8450 1.7000 3.5800 1.7000 3.5800 2.1200 4.0600 2.1200 4.0600 1.7400 4.9650 1.7400
                 4.9650 1.1200 5.0250 1.1200 5.0250 0.6600 5.1450 0.6600 5.1450 1.2400 5.0850 1.2400
                 5.0850 1.6200 5.2450 1.6200 ;
        POLYGON  4.6050 1.1800 3.9400 1.1800 3.9400 2.0000 3.7000 2.0000 3.7000 1.8800 3.8200 1.8800
                 3.8200 0.8800 3.6400 0.8800 3.6400 0.6400 3.7600 0.6400 3.7600 0.7600 3.9400 0.7600
                 3.9400 1.0600 4.6050 1.0600 ;
        POLYGON  3.0000 1.5800 2.6800 1.5800 2.6800 1.4600 2.8800 1.4600 2.8800 0.5200 1.8050 0.5200
                 1.8050 0.6800 1.7700 0.6800 1.7700 0.8000 1.9650 0.8000 1.9650 1.6500 1.7100 1.6500
                 1.7100 1.5300 1.8450 1.5300 1.8450 0.9200 1.6500 0.9200 1.6500 0.5600 1.6850 0.5600
                 1.6850 0.4000 2.3600 0.4000 2.3600 0.3600 2.6000 0.3600 2.6000 0.4000 3.0000 0.4000 ;
        POLYGON  2.2800 2.0600 2.1600 2.0600 2.1600 1.8900 0.8100 1.8900 0.8100 1.6500 0.6450 1.6500
                 0.6450 0.8600 0.5300 0.8600 0.5300 0.7400 0.7700 0.7400 0.7700 0.8600 0.7650 0.8600
                 0.7650 1.5300 0.9300 1.5300 0.9300 1.7700 2.1600 1.7700 2.1600 0.6400 2.2800 0.6400 ;
    END
END SDFFTRX4

MACRO SDFFTRX2
    CLASS CORE ;
    FOREIGN SDFFTRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7100 0.8850 2.8300 1.4400 ;
        RECT  2.6800 0.8850 2.8300 1.2600 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7400 1.1600 7.8850 1.4000 ;
        RECT  7.6100 1.1750 7.7850 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5850 1.1700 9.9650 1.3600 ;
        RECT  9.5850 1.1650 9.8450 1.3800 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1450 1.2300 10.4250 1.4050 ;
        RECT  10.2550 1.0550 10.3900 1.4050 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.6250 0.8550 10.7450 1.2600 ;
        RECT  10.5100 0.5800 10.6600 0.9750 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.8850 1.3800 1.1450 ;
        RECT  1.2300 0.7400 1.3500 2.2100 ;
        RECT  1.0700 0.7400 1.3500 0.8600 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0300 0.7400 2.2700 0.8600 ;
        RECT  2.0700 1.1750 2.2500 1.4350 ;
        RECT  2.0700 0.7400 2.1900 2.2100 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.1250 -0.1800 10.2450 0.9200 ;
        RECT  7.8650 -0.1800 7.9850 0.8400 ;
        RECT  5.7550 -0.1800 5.9950 0.3800 ;
        RECT  3.8750 0.6400 4.1150 0.7600 ;
        RECT  3.9950 -0.1800 4.1150 0.7600 ;
        RECT  2.5100 -0.1800 2.7500 0.3800 ;
        RECT  1.5500 -0.1800 1.7900 0.3800 ;
        RECT  0.6500 -0.1800 0.7700 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.9650 1.6200 11.0850 2.7900 ;
        RECT  10.0650 2.1000 10.1850 2.7900 ;
        RECT  7.7650 1.8400 7.8850 2.7900 ;
        RECT  5.7150 2.2000 5.8350 2.7900 ;
        RECT  3.8750 1.9800 4.1150 2.1000 ;
        RECT  3.8750 1.9800 3.9950 2.7900 ;
        RECT  2.4900 1.5600 2.6100 2.7900 ;
        RECT  1.6500 1.5800 1.7700 2.7900 ;
        RECT  0.8100 1.5600 0.9300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.9850 1.5000 10.6650 1.5000 10.6650 1.9800 8.8250 1.9800 8.8250 1.7200 9.1050 1.7200
                 9.1050 0.8400 8.9850 0.8400 8.9850 0.6000 9.1050 0.6000 9.1050 0.7200 9.2250 0.7200
                 9.2250 1.8600 10.5450 1.8600 10.5450 1.3800 10.8650 1.3800 10.8650 0.6800
                 10.9850 0.6800 ;
        POLYGON  9.8250 0.9200 9.4650 0.9200 9.4650 1.5000 9.7050 1.5000 9.7050 1.7400 9.5850 1.7400
                 9.5850 1.6200 9.3450 1.6200 9.3450 0.8000 9.7050 0.8000 9.7050 0.6800 9.3450 0.6800
                 9.3450 0.4800 8.8650 0.4800 8.8650 0.9800 8.9850 0.9800 8.9850 1.1000 8.8650 1.1000
                 8.8650 1.3200 8.3650 1.3200 8.3650 1.4800 8.2450 1.4800 8.2450 1.2000 8.7450 1.2000
                 8.7450 0.3600 9.4650 0.3600 9.4650 0.5600 9.8250 0.5600 ;
        POLYGON  8.6250 1.0800 8.1250 1.0800 8.1250 1.6000 8.5250 1.6000 8.5250 1.9600 8.4050 1.9600
                 8.4050 1.7200 7.1750 1.7200 7.1750 1.7800 6.8950 1.7800 6.8950 1.6600 7.0550 1.6600
                 7.0550 0.6800 7.1750 0.6800 7.1750 1.6000 8.0050 1.6000 8.0050 0.9600 8.5050 0.9600
                 8.5050 0.6000 8.6250 0.6000 ;
        POLYGON  7.5650 0.8400 7.4450 0.8400 7.4450 0.6000 7.3450 0.6000 7.3450 0.5600 6.9350 0.5600
                 6.9350 1.1000 6.7750 1.1000 6.7750 1.2800 6.9350 1.2800 6.9350 1.5200 6.7750 1.5200
                 6.7750 1.9000 7.5250 1.9000 7.5250 2.0200 6.6550 2.0200 6.6550 0.9800 6.8150 0.9800
                 6.8150 0.5600 6.2900 0.5600 6.2900 0.6200 5.1550 0.6200 5.1550 1.2600 5.0350 1.2600
                 5.0350 0.5000 6.1700 0.5000 6.1700 0.4400 6.3150 0.4400 6.3150 0.4200 6.5550 0.4200
                 6.5550 0.4400 7.4650 0.4400 7.4650 0.4800 7.5650 0.4800 ;
        POLYGON  6.6950 0.8600 6.5350 0.8600 6.5350 1.8400 6.4150 1.8400 6.4150 1.4400 5.5350 1.4400
                 5.5350 1.3200 6.4150 1.3200 6.4150 0.7400 6.6950 0.7400 ;
        POLYGON  6.4550 2.2200 6.1450 2.2200 6.1450 2.0800 5.2750 2.0800 5.2750 2.2200 5.0350 2.2200
                 5.0350 2.0800 4.5550 2.0800 4.5550 1.8600 2.9700 1.8600 2.9700 0.7400 3.2300 0.7400
                 3.2300 0.8600 3.0900 0.8600 3.0900 1.7400 4.5550 1.7400 4.5550 1.2400 4.4350 1.2400
                 4.4350 1.1200 4.6750 1.1200 4.6750 1.9600 6.2650 1.9600 6.2650 2.1000 6.4550 2.1000 ;
        POLYGON  6.1150 1.2000 5.4150 1.2000 5.4150 1.7200 5.3550 1.7200 5.3550 1.8400 5.2350 1.8400
                 5.2350 1.6000 5.2950 1.6000 5.2950 0.8600 5.2750 0.8600 5.2750 0.7400 5.5150 0.7400
                 5.5150 0.8600 5.4150 0.8600 5.4150 1.0800 6.1150 1.0800 ;
        POLYGON  4.9350 1.8400 4.8150 1.8400 4.8150 1.5000 4.7950 1.5000 4.7950 0.9200 4.4250 0.9200
                 4.4250 1.0000 3.8950 1.0000 3.8950 1.2600 3.7750 1.2600 3.7750 0.8800 4.3050 0.8800
                 4.3050 0.8000 4.7750 0.8000 4.7750 0.6800 4.8950 0.6800 4.8950 0.8000 4.9150 0.8000
                 4.9150 1.3800 4.9350 1.3800 ;
        POLYGON  4.3150 1.4400 4.1350 1.4400 4.1350 1.5000 3.6350 1.5000 3.6350 1.6200 3.3950 1.6200
                 3.3950 1.5000 3.5150 1.5000 3.5150 0.6200 2.5100 0.6200 2.5100 1.2400 2.3700 1.2400
                 2.3700 1.0000 2.3900 1.0000 2.3900 0.6200 1.9100 0.6200 1.9100 1.4600 1.7900 1.4600
                 1.7900 0.6200 0.3900 0.6200 0.3900 0.5200 0.2700 0.5200 0.2700 0.4000 0.5100 0.4000
                 0.5100 0.5000 3.6350 0.5000 3.6350 1.3800 4.0150 1.3800 4.0150 1.3200 4.3150 1.3200 ;
        POLYGON  1.1100 1.1800 0.4500 1.1800 0.4500 1.8000 0.3300 1.8000 0.3300 0.8600 0.1100 0.8600
                 0.1100 0.7400 0.4500 0.7400 0.4500 1.0600 1.1100 1.0600 ;
    END
END SDFFTRX2

MACRO SDFFTRX1
    CLASS CORE ;
    FOREIGN SDFFTRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0050 1.2200 2.1250 1.4600 ;
        RECT  1.7550 1.5200 2.0150 1.6700 ;
        RECT  1.8950 1.3400 2.0150 1.6700 ;
        END
    END CK
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7400 1.1850 7.0150 1.4350 ;
        RECT  6.7400 1.1650 6.8900 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7150 0.9400 8.9750 1.0900 ;
        RECT  8.7150 0.9400 8.9550 1.3000 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 1.1650 9.5550 1.3800 ;
        RECT  9.2150 0.9800 9.3350 1.3600 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.7750 0.8850 10.0800 1.2200 ;
        RECT  9.9300 0.8800 10.0800 1.2200 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 2.2100 ;
        RECT  1.2300 0.8850 1.4850 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  9.0750 -0.1800 9.1950 0.8200 ;
        RECT  6.9950 -0.1800 7.1150 0.8400 ;
        RECT  4.8850 -0.1800 5.1250 0.3200 ;
        RECT  3.1050 -0.1800 3.3450 0.3200 ;
        RECT  1.7850 -0.1800 1.9050 0.7300 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  9.9150 1.5800 10.0350 2.7900 ;
        RECT  9.0150 2.0600 9.1350 2.7900 ;
        RECT  6.9950 1.8800 7.1150 2.7900 ;
        RECT  4.9450 2.1400 5.0650 2.7900 ;
        RECT  3.2850 2.0800 3.5250 2.2000 ;
        RECT  3.2850 2.0800 3.4050 2.7900 ;
        RECT  1.7850 1.7900 1.9050 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.3200 1.4600 9.7950 1.4600 9.7950 1.6200 9.6150 1.6200 9.6150 1.8600 9.2350 1.8600
                 9.2350 1.9400 8.1750 1.9400 8.1750 2.0000 8.0550 2.0000 8.0550 1.4400 8.2350 1.4400
                 8.2350 0.8400 8.1150 0.8400 8.1150 0.6000 8.2350 0.6000 8.2350 0.7200 8.3550 0.7200
                 8.3550 1.5600 8.1750 1.5600 8.1750 1.8200 9.1150 1.8200 9.1150 1.7400 9.4950 1.7400
                 9.4950 1.5000 9.6750 1.5000 9.6750 1.3400 10.2000 1.3400 10.2000 0.7600 9.6550 0.7600
                 9.6550 0.6400 10.3200 0.6400 ;
        POLYGON  8.7750 0.8200 8.5950 0.8200 8.5950 1.4200 8.6550 1.4200 8.6550 1.7000 8.5350 1.7000
                 8.5350 1.5400 8.4750 1.5400 8.4750 0.7000 8.6550 0.7000 8.6550 0.4800 7.9950 0.4800
                 7.9950 0.9800 8.1150 0.9800 8.1150 1.1000 7.9950 1.1000 7.9950 1.3200 7.4950 1.3200
                 7.4950 1.4400 7.3750 1.4400 7.3750 1.2000 7.8750 1.2000 7.8750 0.3600 8.7750 0.3600 ;
        POLYGON  7.7550 1.0800 7.2550 1.0800 7.2550 1.5600 7.7550 1.5600 7.7550 2.0000 7.6350 2.0000
                 7.6350 1.6800 6.3650 1.6800 6.3650 1.7200 6.1250 1.7200 6.1250 1.6000 6.2450 1.6000
                 6.2450 0.9200 6.1850 0.9200 6.1850 0.6800 6.3050 0.6800 6.3050 0.8000 6.3650 0.8000
                 6.3650 1.5600 7.1350 1.5600 7.1350 0.9600 7.6350 0.9600 7.6350 0.6000 7.7550 0.6000 ;
        POLYGON  6.7550 1.9600 5.8850 1.9600 5.8850 0.9800 5.9450 0.9800 5.9450 0.5600 4.3450 0.5600
                 4.3450 1.2400 4.2250 1.2400 4.2250 0.4400 5.4250 0.4400 5.4250 0.4000 5.6650 0.4000
                 5.6650 0.4400 6.5450 0.4400 6.5450 0.4800 6.6950 0.4800 6.6950 0.8400 6.5750 0.8400
                 6.5750 0.6000 6.4250 0.6000 6.4250 0.5600 6.0650 0.5600 6.0650 1.1000 6.0050 1.1000
                 6.0050 1.2800 6.1250 1.2800 6.1250 1.4000 6.0050 1.4000 6.0050 1.8400 6.7550 1.8400 ;
        POLYGON  5.8250 0.8600 5.7650 0.8600 5.7650 1.7800 5.6450 1.7800 5.6450 1.4400 4.8250 1.4400
                 4.8250 1.4000 4.7050 1.4000 4.7050 1.2800 4.9450 1.2800 4.9450 1.3200 5.6450 1.3200
                 5.6450 0.8600 5.5850 0.8600 5.5850 0.7400 5.8250 0.7400 ;
        POLYGON  5.6850 2.1600 5.4450 2.1600 5.4450 2.0200 4.3650 2.0200 4.3650 2.1600 4.1250 2.1600
                 4.1250 2.0200 3.6450 2.0200 3.6450 1.9600 2.5300 1.9600 2.5300 1.9200 2.2650 1.9200
                 2.2650 0.6800 2.3850 0.6800 2.3850 1.8000 2.6500 1.8000 2.6500 1.8400 3.6450 1.8400
                 3.6450 1.1800 3.6250 1.1800 3.6250 1.0600 3.8650 1.0600 3.8650 1.1800 3.7650 1.1800
                 3.7650 1.9000 5.5650 1.9000 5.5650 2.0400 5.6850 2.0400 ;
        POLYGON  5.3450 1.2000 5.1050 1.2000 5.1050 1.1600 4.5850 1.1600 4.5850 1.7800 4.4650 1.7800
                 4.4650 0.6800 4.5850 0.6800 4.5850 1.0400 5.2250 1.0400 5.2250 1.0800 5.3450 1.0800 ;
        POLYGON  4.1650 1.7800 4.0450 1.7800 4.0450 1.4800 3.9850 1.4800 3.9850 0.9200 3.8250 0.9200
                 3.8250 0.6800 2.8950 0.6800 2.8950 0.5600 2.7450 0.5600 2.7450 0.4000 2.9850 0.4000
                 2.9850 0.4400 3.0150 0.4400 3.0150 0.5600 3.9450 0.5600 3.9450 0.8000 4.1050 0.8000
                 4.1050 1.3600 4.1650 1.3600 ;
        POLYGON  3.5050 1.1800 2.9250 1.1800 2.9250 1.6000 3.0450 1.6000 3.0450 1.7200 2.8050 1.7200
                 2.8050 0.9200 2.6550 0.9200 2.6550 0.8000 2.5050 0.8000 2.5050 0.5600 2.1450 0.5600
                 2.1450 0.9700 1.7650 0.9700 1.7650 1.2400 1.6450 1.2400 1.6450 0.8500 2.0250 0.8500
                 2.0250 0.4400 2.6250 0.4400 2.6250 0.6800 2.7750 0.6800 2.7750 0.8000 2.9250 0.8000
                 2.9250 1.0600 3.5050 1.0600 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END SDFFTRX1

MACRO SDFFSXL
    CLASS CORE ;
    FOREIGN SDFFSXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5850 0.3600 5.7050 0.6000 ;
        RECT  4.8400 0.4600 5.7050 0.5800 ;
        RECT  3.7800 0.4200 4.9600 0.4800 ;
        RECT  4.5750 0.4600 5.7050 0.5400 ;
        RECT  3.7800 0.3600 4.6950 0.4800 ;
        RECT  3.7800 0.3600 3.9000 1.3400 ;
        RECT  3.6350 1.2200 3.9000 1.3400 ;
        RECT  3.4950 1.2300 3.7550 1.3800 ;
        RECT  3.0800 1.2300 3.7550 1.3500 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2750 0.9700 8.5950 1.1150 ;
        RECT  8.1350 0.9100 8.3950 1.0900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7150 0.8700 8.9750 1.1000 ;
        RECT  8.7550 0.8700 8.8750 1.2800 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.0750 1.2100 10.1950 1.6200 ;
        RECT  9.8750 1.2300 10.1950 1.4600 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3950 0.9700 10.5950 1.0900 ;
        RECT  10.1650 0.9400 10.4250 1.0900 ;
        RECT  9.8350 0.8700 9.9550 1.1100 ;
        RECT  9.2350 1.4900 9.5150 1.6100 ;
        RECT  9.3950 0.9700 9.5150 1.6100 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1644  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8150 0.8850 1.0900 1.1450 ;
        RECT  0.8150 0.7400 0.9950 1.1450 ;
        RECT  0.8150 0.7400 0.9350 2.1350 ;
        RECT  0.7550 0.7400 0.9950 0.8600 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1644  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9900 0.7400 2.2300 0.8600 ;
        RECT  1.9900 0.7400 2.1100 1.5050 ;
        RECT  1.8100 1.4650 2.0150 1.6250 ;
        RECT  1.8400 1.3850 2.1100 1.5050 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.3150 -0.1800 10.4350 0.7500 ;
        RECT  8.7550 -0.1800 8.8750 0.7500 ;
        RECT  6.5650 -0.1800 6.6850 0.6500 ;
        RECT  5.1850 -0.1800 5.4250 0.3400 ;
        RECT  2.9200 -0.1800 3.0400 0.7100 ;
        RECT  1.5100 -0.1800 1.6300 0.4000 ;
        RECT  0.1550 0.7400 0.3950 0.8600 ;
        RECT  0.1550 -0.1800 0.2750 0.8600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.1950 1.9800 10.3150 2.7900 ;
        RECT  8.7550 1.9700 8.8750 2.7900 ;
        RECT  6.6650 2.1100 6.7850 2.7900 ;
        RECT  5.6450 2.2900 5.8850 2.7900 ;
        RECT  3.3950 2.0300 3.6350 2.1500 ;
        RECT  3.3950 2.0300 3.5150 2.7900 ;
        RECT  2.6150 1.9700 2.7350 2.7900 ;
        RECT  1.4750 1.5050 1.5950 2.7900 ;
        RECT  0.3950 1.9700 0.5150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.8550 0.7500 10.8350 0.7500 10.8350 1.9700 10.7950 1.9700 10.7950 2.0900
                 10.6750 2.0900 10.6750 1.8600 9.6350 1.8600 9.6350 1.5300 9.7550 1.5300 9.7550 1.7400
                 10.7150 1.7400 10.7150 0.6300 10.7350 0.6300 10.7350 0.5100 10.8550 0.5100 ;
        POLYGON  9.7950 0.7500 9.2750 0.7500 9.2750 1.3700 9.1150 1.3700 9.1150 1.7300 9.5150 1.7300
                 9.5150 2.0900 9.3950 2.0900 9.3950 1.8500 7.8950 1.8500 7.8950 1.6900 7.8450 1.6900
                 7.8450 1.5700 7.8950 1.5700 7.8950 0.7200 7.8250 0.7200 7.8250 0.6000 8.0650 0.6000
                 8.0650 0.7200 8.0150 0.7200 8.0150 1.5700 8.0850 1.5700 8.0850 1.7300 8.9950 1.7300
                 8.9950 1.2500 9.1550 1.2500 9.1550 0.6300 9.6750 0.6300 9.6750 0.5100 9.7950 0.5100 ;
        POLYGON  8.5150 2.0900 7.3250 2.0900 7.3250 2.2100 7.2050 2.2100 7.2050 2.0900 7.0350 2.0900
                 7.0350 1.9900 6.3600 1.9900 6.3600 2.1700 5.3250 2.1700 5.3250 2.0500 6.2400 2.0500
                 6.2400 1.8700 7.1550 1.8700 7.1550 1.9700 7.6050 1.9700 7.6050 1.1200 7.5850 1.1200
                 7.5850 0.3600 8.3950 0.3600 8.3950 0.7500 8.2750 0.7500 8.2750 0.4800 7.7050 0.4800
                 7.7050 0.8800 7.7650 0.8800 7.7650 1.1200 7.7250 1.1200 7.7250 1.9700 8.5150 1.9700 ;
        POLYGON  7.4850 1.7500 7.3650 1.7500 7.3650 1.3700 6.3850 1.3700 6.3850 1.2500 7.3450 1.2500
                 7.3450 0.5400 7.4650 0.5400 7.4650 1.2500 7.4850 1.2500 ;
        POLYGON  7.2250 1.1200 7.1050 1.1200 7.1050 0.8900 6.3250 0.8900 6.3250 0.5600 5.9450 0.5600
                 5.9450 1.0200 5.4050 1.0200 5.4050 1.6900 5.1650 1.6900 5.1650 1.5700 5.2850 1.5700
                 5.2850 1.0200 4.6200 1.0200 4.6200 1.1600 4.5000 1.1600 4.5000 0.9000 4.7800 0.9000
                 4.7800 0.7400 5.0200 0.7400 5.0200 0.9000 5.8250 0.9000 5.8250 0.4400 6.4450 0.4400
                 6.4450 0.7700 7.2250 0.7700 ;
        POLYGON  6.9650 1.1300 6.2050 1.1300 6.2050 1.5100 6.3050 1.5100 6.3050 1.7500 5.7750 1.7500
                 5.7750 1.9300 4.8350 1.9300 4.8350 1.4000 4.2600 1.4000 4.2600 0.6600 4.6200 0.6600
                 4.6200 0.7800 4.3800 0.7800 4.3800 1.2800 4.9550 1.2800 4.9550 1.8100 5.6550 1.8100
                 5.6550 1.6300 6.0850 1.6300 6.0850 0.6800 6.2050 0.6800 6.2050 1.0100 6.9650 1.0100 ;
        POLYGON  4.5350 1.8200 4.4150 1.8200 4.4150 1.6400 2.7000 1.6400 2.7000 1.0700 2.8200 1.0700
                 2.8200 1.5200 4.0200 1.5200 4.0200 0.6000 4.1400 0.6000 4.1400 1.5200 4.5350 1.5200 ;
        POLYGON  4.1750 1.8800 4.0550 1.8800 4.0550 1.9100 3.2600 1.9100 3.2600 2.0300 2.9750 2.0300
                 2.9750 1.9100 3.1400 1.9100 3.1400 1.7900 3.9350 1.7900 3.9350 1.7600 4.1750 1.7600 ;
        POLYGON  3.6600 1.1000 3.4200 1.1000 3.4200 0.9500 2.5600 0.9500 2.5600 1.8500 2.3750 1.8500
                 2.3750 2.0750 2.1350 2.0750 2.1350 1.7300 2.4400 1.7300 2.4400 0.6200 1.8700 0.6200
                 1.8700 1.1800 1.6300 1.1800 1.6300 1.0600 1.7500 1.0600 1.7500 0.5000 2.5600 0.5000
                 2.5600 0.8300 3.5400 0.8300 3.5400 0.9800 3.6600 0.9800 ;
        POLYGON  1.3300 1.3850 1.1750 1.3850 1.1750 1.6250 1.0550 1.6250 1.0550 1.2650 1.2100 1.2650
                 1.2100 0.6200 0.6350 0.6200 0.6350 1.0000 0.6550 1.0000 0.6550 1.2400 0.5150 1.2400
                 0.5150 0.5000 1.3300 0.5000 ;
    END
END SDFFSXL

MACRO SDFFSX4
    CLASS CORE ;
    FOREIGN SDFFSX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.2100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4200 0.5900 1.5400 2.2100 ;
        RECT  0.5800 1.3150 1.5400 1.4350 ;
        RECT  0.5800 1.1750 0.8000 1.4350 ;
        RECT  0.5800 0.5900 0.7000 2.2100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8900 0.6800 4.0100 2.1400 ;
        RECT  2.9700 1.0250 4.0100 1.1450 ;
        RECT  3.0500 0.6800 3.1700 2.1400 ;
        RECT  2.9700 0.8850 3.1700 1.1450 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1650 0.5200 8.2850 0.9800 ;
        RECT  7.4600 0.5200 8.2850 0.6400 ;
        RECT  7.4600 0.3600 7.5800 0.6400 ;
        RECT  5.8700 0.3600 7.5800 0.4800 ;
        RECT  5.8700 0.8850 6.0200 1.1450 ;
        RECT  5.2500 1.2400 5.9900 1.3600 ;
        RECT  5.8700 0.3600 5.9900 1.3600 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.1750 1.5000 11.5650 1.6200 ;
        RECT  11.0350 1.5200 11.2950 1.6700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.7250 1.2600 11.8450 1.5000 ;
        RECT  11.3250 1.2600 11.8450 1.3800 ;
        RECT  11.3250 1.2300 11.5850 1.3800 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.0650 1.2300 13.3250 1.5000 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.7000 1.1750 13.8500 1.4350 ;
        RECT  13.5250 1.1700 13.8200 1.2900 ;
        RECT  13.5250 0.9900 13.6450 1.2900 ;
        RECT  12.4050 0.9900 13.6450 1.1100 ;
        RECT  12.7050 0.9900 12.9450 1.1300 ;
        RECT  12.2050 1.4400 12.5250 1.5600 ;
        RECT  12.4050 0.9900 12.5250 1.5600 ;
        RECT  12.2050 1.4400 12.3250 1.6800 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.2100 0.1800 ;
        RECT  13.2650 -0.1800 13.3850 0.8700 ;
        RECT  11.9250 -0.1800 12.0450 0.6300 ;
        RECT  11.0250 -0.1800 11.2650 0.3300 ;
        RECT  9.0350 -0.1800 9.1550 0.8500 ;
        RECT  7.8850 -0.1800 8.1250 0.4000 ;
        RECT  5.0900 0.6000 5.3300 0.7200 ;
        RECT  5.2100 -0.1800 5.3300 0.7200 ;
        RECT  4.3100 -0.1800 4.4300 0.7800 ;
        RECT  3.4700 -0.1800 3.5900 0.7300 ;
        RECT  2.6300 -0.1800 2.7500 0.7300 ;
        RECT  1.9000 -0.1800 2.0200 0.5300 ;
        RECT  1.0000 -0.1800 1.1200 0.6400 ;
        RECT  0.1600 -0.1800 0.2800 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.2100 2.7900 ;
        RECT  13.1850 1.9000 13.3050 2.7900 ;
        RECT  11.7250 1.9000 11.8450 2.7900 ;
        RECT  10.9150 2.1700 11.0350 2.7900 ;
        RECT  8.7450 2.2900 8.9850 2.7900 ;
        RECT  7.5450 2.1200 7.7850 2.2400 ;
        RECT  7.5450 2.1200 7.6650 2.7900 ;
        RECT  5.9900 1.9600 6.2300 2.0800 ;
        RECT  5.9900 1.9600 6.1100 2.7900 ;
        RECT  5.1500 1.7200 5.2700 2.7900 ;
        RECT  4.3100 1.6200 4.4300 2.7900 ;
        RECT  3.4700 1.4900 3.5900 2.7900 ;
        RECT  2.6300 1.4900 2.7500 2.7900 ;
        RECT  1.8400 1.9700 1.9600 2.7900 ;
        RECT  1.0000 1.5600 1.1200 2.7900 ;
        RECT  0.1600 1.5600 0.2800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.0900 1.8600 13.7250 1.8600 13.7250 2.0200 13.6050 2.0200 13.6050 1.7400
                 12.6450 1.7400 12.6450 1.4600 12.7650 1.4600 12.7650 1.6200 13.9700 1.6200
                 13.9700 0.8100 13.6250 0.8100 13.6250 0.6900 14.0900 0.6900 ;
        POLYGON  12.8050 0.8100 12.3500 0.8100 12.3500 0.8700 12.0850 0.8700 12.0850 1.8000
                 12.4850 1.8000 12.4850 2.0400 12.3650 2.0400 12.3650 1.9200 11.9650 1.9200
                 11.9650 0.8700 11.6850 0.8700 11.6850 0.5700 10.7850 0.5700 10.7850 0.4800
                 10.2150 0.4800 10.2150 1.2100 10.1650 1.2100 10.1650 1.7500 10.0450 1.7500
                 10.0450 1.0900 10.0950 1.0900 10.0950 0.3600 10.9050 0.3600 10.9050 0.4500
                 11.8050 0.4500 11.8050 0.7500 12.2300 0.7500 12.2300 0.6900 12.8050 0.6900 ;
        POLYGON  11.5650 0.8100 11.4450 0.8100 11.4450 0.9800 10.8350 0.9800 10.8350 1.1000
                 10.7950 1.1000 10.7950 1.8400 11.4050 1.8400 11.4050 1.9600 10.7950 1.9600
                 10.7950 2.2500 10.0800 2.2500 10.0800 2.2300 9.5500 2.2300 9.5500 2.1700 7.9050 2.1700
                 7.9050 2.0000 6.7400 2.0000 6.7400 1.4000 6.3800 1.4000 6.3800 1.0800 6.5000 1.0800
                 6.5000 1.2800 6.8600 1.2800 6.8600 1.8800 8.0250 1.8800 8.0250 2.0500 9.6700 2.0500
                 9.6700 2.1100 10.2000 2.1100 10.2000 2.1300 10.6750 2.1300 10.6750 0.8600
                 11.3250 0.8600 11.3250 0.6900 11.5650 0.6900 ;
        POLYGON  10.6650 0.7200 10.5550 0.7200 10.5550 2.0100 10.4350 2.0100 10.4350 1.9900
                 9.8050 1.9900 9.8050 1.9300 8.1450 1.9300 8.1450 1.7600 7.3000 1.7600 7.3000 1.2400
                 7.2200 1.2400 7.2200 1.0000 7.3400 1.0000 7.3400 1.1200 7.4200 1.1200 7.4200 1.6400
                 8.2650 1.6400 8.2650 1.8100 9.8050 1.8100 9.8050 1.4500 9.7650 1.4500 9.7650 1.1700
                 9.8850 1.1700 9.8850 1.3300 9.9250 1.3300 9.9250 1.8700 10.4350 1.8700 10.4350 0.7200
                 10.4250 0.7200 10.4250 0.6000 10.6650 0.6000 ;
        POLYGON  9.7950 0.8500 9.5650 0.8500 9.5650 1.5700 9.6850 1.5700 9.6850 1.6900 9.4450 1.6900
                 9.4450 1.3500 8.6450 1.3500 8.6450 1.2300 9.4450 1.2300 9.4450 0.7300 9.6750 0.7300
                 9.6750 0.6100 9.7950 0.6100 ;
        POLYGON  9.2250 1.1100 8.5250 1.1100 8.5250 1.5700 8.6250 1.5700 8.6250 1.6900 8.3850 1.6900
                 8.3850 1.5700 8.4050 1.5700 8.4050 1.2200 7.7600 1.2200 7.7600 1.4000 7.8800 1.4000
                 7.8800 1.5200 7.6400 1.5200 7.6400 0.8800 6.9400 0.8800 6.9400 0.7200 6.8200 0.7200
                 6.8200 0.6000 7.0600 0.6000 7.0600 0.7600 7.7600 0.7600 7.7600 1.1000 8.4050 1.1000
                 8.4050 0.9900 8.6450 0.9900 8.6450 0.4000 8.7650 0.4000 8.7650 0.9900 9.2250 0.9900 ;
        POLYGON  7.1800 1.6000 7.0600 1.6000 7.0600 1.4800 6.9800 1.4800 6.9800 1.1600 6.7000 1.1600
                 6.7000 0.9600 6.2600 0.9600 6.2600 1.6000 5.0100 1.6000 5.0100 1.5400 4.9700 1.5400
                 4.9700 1.3000 5.0900 1.3000 5.0900 1.4200 5.1300 1.4200 5.1300 1.4800 6.1400 1.4800
                 6.1400 0.8400 6.4000 0.8400 6.4000 0.6000 6.6400 0.6000 6.6400 0.7200 6.5200 0.7200
                 6.5200 0.8400 6.8200 0.8400 6.8200 1.0400 7.1000 1.0400 7.1000 1.3600 7.1800 1.3600 ;
        POLYGON  6.6200 1.6400 6.5000 1.6400 6.5000 1.8400 5.8100 1.8400 5.8100 1.9600 5.5700 1.9600
                 5.5700 1.8400 5.6900 1.8400 5.6900 1.7200 6.3800 1.7200 6.3800 1.5200 6.6200 1.5200 ;
        POLYGON  5.7500 1.1200 4.8500 1.1200 4.8500 2.1400 4.7300 2.1400 4.7300 1.1200 4.2900 1.1200
                 4.2900 1.2400 4.1700 1.2400 4.1700 1.0000 4.7300 1.0000 4.7300 0.6400 4.8500 0.6400
                 4.8500 1.0000 5.6300 1.0000 5.6300 0.8800 5.7500 0.8800 ;
        POLYGON  2.3300 1.8200 2.2100 1.8200 2.2100 1.4200 1.6600 1.4200 1.6600 1.3000 2.2100 1.3000
                 2.2100 0.6800 2.3300 0.6800 ;
    END
END SDFFSX4

MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.2750 0.3600 6.5150 0.4800 ;
        RECT  5.6950 0.8500 6.4150 0.9700 ;
        RECT  6.2950 0.3600 6.4150 0.9700 ;
        RECT  5.6950 0.3800 5.8150 0.9700 ;
        RECT  4.3650 0.3600 5.8100 0.4800 ;
        RECT  5.6900 0.3800 5.8150 0.5000 ;
        RECT  4.3650 1.2300 4.6250 1.3800 ;
        RECT  4.3650 0.3600 4.4850 1.3800 ;
        RECT  3.6850 1.2400 4.6250 1.3600 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.1450 0.8450 9.4650 1.0100 ;
        RECT  9.0050 0.8900 9.2650 1.0900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5850 0.7750 9.8250 0.9800 ;
        RECT  9.6400 0.7600 9.7900 1.1550 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7850 1.2600 11.2950 1.3850 ;
        RECT  11.0350 1.2300 11.2950 1.3850 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1850 0.9250 11.2250 1.0450 ;
        RECT  10.7450 0.9250 11.0050 1.0900 ;
        RECT  10.4450 0.7600 10.5650 1.0450 ;
        RECT  10.0650 1.5150 10.3050 1.6350 ;
        RECT  10.1850 0.9250 10.3050 1.6350 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.5900 0.6750 2.2100 ;
        RECT  0.3600 0.8850 0.6750 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1950 0.6800 2.3150 1.9900 ;
        RECT  2.1000 1.1750 2.3150 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  10.9250 -0.1800 11.0450 0.6400 ;
        RECT  9.6450 -0.1800 9.7650 0.6400 ;
        RECT  7.3550 -0.1800 7.4750 0.5800 ;
        RECT  5.9350 0.6100 6.1750 0.7300 ;
        RECT  6.0350 -0.1800 6.1550 0.7300 ;
        RECT  3.5250 0.6600 3.7650 0.7800 ;
        RECT  3.5250 -0.1800 3.6450 0.7800 ;
        RECT  2.6150 -0.1800 2.7350 0.7800 ;
        RECT  1.7750 -0.1800 1.8950 0.7300 ;
        RECT  1.0350 -0.1800 1.1550 0.5300 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  10.9250 1.9350 11.0450 2.7900 ;
        RECT  9.5850 1.9950 9.8250 2.1150 ;
        RECT  9.5850 1.9950 9.7050 2.7900 ;
        RECT  7.4550 1.6600 7.5750 2.7900 ;
        RECT  6.4350 2.2900 6.6750 2.7900 ;
        RECT  4.1850 2.0500 4.4250 2.1700 ;
        RECT  4.1850 2.0500 4.3050 2.7900 ;
        RECT  3.3450 1.9700 3.4650 2.7900 ;
        RECT  2.6750 2.1400 2.7950 2.7900 ;
        RECT  1.7150 1.9800 1.8350 2.7900 ;
        RECT  0.9750 1.7300 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.5350 1.7450 11.4650 1.7450 11.4650 2.0550 11.3450 2.0550 11.3450 1.6250
                 10.5450 1.6250 10.5450 1.3750 10.4250 1.3750 10.4250 1.2550 10.6650 1.2550
                 10.6650 1.5050 11.4150 1.5050 11.4150 1.1100 11.3450 1.1100 11.3450 0.4000
                 11.4650 0.4000 11.4650 0.9900 11.5350 0.9900 ;
        POLYGON  10.4050 0.6400 10.0650 0.6400 10.0650 1.3950 9.9450 1.3950 9.9450 1.7550
                 10.4050 1.7550 10.4050 2.0550 10.2850 2.0550 10.2850 1.8750 8.7550 1.8750
                 8.7550 1.7600 8.6350 1.7600 8.6350 1.6400 8.7550 1.6400 8.7550 0.7200 8.6950 0.7200
                 8.6950 0.6000 8.9350 0.6000 8.9350 0.7200 8.8750 0.7200 8.8750 1.7550 9.8250 1.7550
                 9.8250 1.2750 9.9450 1.2750 9.9450 0.5200 10.2850 0.5200 10.2850 0.4000 10.4050 0.4000 ;
        POLYGON  9.4050 2.1150 8.3950 2.1150 8.3950 1.9900 8.1750 1.9900 8.1750 2.1500 7.9350 2.1500
                 7.9350 1.9900 7.7450 1.9900 7.7450 1.5400 7.3350 1.5400 7.3350 2.1100 6.8050 2.1100
                 6.8050 2.1700 6.1150 2.1700 6.1150 2.0500 6.6850 2.0500 6.6850 1.9900 7.2150 1.9900
                 7.2150 1.4200 7.8650 1.4200 7.8650 1.8700 8.3950 1.8700 8.3950 1.4000 8.4550 1.4000
                 8.4550 0.3600 9.2650 0.3600 9.2650 0.6400 9.1450 0.6400 9.1450 0.4800 8.5750 0.4800
                 8.5750 1.5200 8.5150 1.5200 8.5150 1.9950 9.4050 1.9950 ;
        POLYGON  8.3350 1.2800 8.2750 1.2800 8.2750 1.7500 8.1550 1.7500 8.1550 1.3000 7.1750 1.3000
                 7.1750 1.1800 8.1550 1.1800 8.1550 1.1600 8.2150 1.1600 8.2150 0.7200 8.0950 0.7200
                 8.0950 0.6000 8.3350 0.6000 ;
        POLYGON  8.0950 1.0400 7.8550 1.0400 7.8550 0.8200 7.1150 0.8200 7.1150 0.5000 6.7550 0.5000
                 6.7550 0.7200 6.6550 0.7200 6.6550 1.2100 6.0750 1.2100 6.0750 1.5700 6.1950 1.5700
                 6.1950 1.6900 5.9550 1.6900 5.9550 1.2100 5.2250 1.2100 5.2250 1.0300 5.4550 1.0300
                 5.4550 0.6200 5.5750 0.6200 5.5750 1.0900 6.5350 1.0900 6.5350 0.6000 6.6350 0.6000
                 6.6350 0.3800 7.2350 0.3800 7.2350 0.7000 7.9750 0.7000 7.9750 0.9200 8.0950 0.9200 ;
        POLYGON  7.7350 1.0600 6.9950 1.0600 6.9950 1.5100 7.0950 1.5100 7.0950 1.8700 6.5650 1.8700
                 6.5650 1.9300 5.6250 1.9300 5.6250 1.4500 4.9850 1.4500 4.9850 0.7200 5.0250 0.7200
                 5.0250 0.6000 5.1450 0.6000 5.1450 0.8400 5.1050 0.8400 5.1050 1.3300 5.7450 1.3300
                 5.7450 1.8100 6.4450 1.8100 6.4450 1.7500 6.9750 1.7500 6.9750 1.6300 6.8750 1.6300
                 6.8750 0.6200 6.9950 0.6200 6.9950 0.9400 7.7350 0.9400 ;
        POLYGON  5.3250 1.8700 5.2050 1.8700 5.2050 1.6900 3.4450 1.6900 3.4450 1.3800 3.2750 1.3800
                 3.2750 1.1400 3.3950 1.1400 3.3950 1.2600 3.5650 1.2600 3.5650 1.5700 4.7450 1.5700
                 4.7450 1.1100 4.6050 1.1100 4.6050 0.6000 4.7250 0.6000 4.7250 0.9900 4.8650 0.9900
                 4.8650 1.5700 5.3250 1.5700 ;
        POLYGON  4.9650 1.9300 3.9450 1.9300 3.9450 2.0300 3.7050 2.0300 3.7050 1.9100 3.8250 1.9100
                 3.8250 1.8100 4.9650 1.8100 ;
        POLYGON  4.2450 1.1200 4.0050 1.1200 4.0050 1.0200 3.1550 1.0200 3.1550 1.8200 3.0350 1.8200
                 3.0350 1.0200 2.5950 1.0200 2.5950 1.2400 2.4750 1.2400 2.4750 0.9000 3.0350 0.9000
                 3.0350 0.6400 3.1550 0.6400 3.1550 0.9000 4.1250 0.9000 4.1250 1.0000 4.2450 1.0000 ;
        POLYGON  1.4150 1.0500 1.4050 1.0500 1.4050 1.5800 1.2850 1.5800 1.2850 1.1700 0.7950 1.1700
                 0.7950 1.0500 1.2850 1.0500 1.2850 0.9300 1.2950 0.9300 1.2950 0.6800 1.4150 0.6800 ;
    END
END SDFFSX2

MACRO SDFFSX1
    CLASS CORE ;
    FOREIGN SDFFSX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7200 0.3600 5.9600 0.4800 ;
        RECT  5.1200 0.8300 5.8400 0.9500 ;
        RECT  5.7200 0.3600 5.8400 0.9500 ;
        RECT  5.1200 0.3800 5.2400 0.9500 ;
        RECT  3.7450 0.3800 5.2400 0.5000 ;
        RECT  3.7450 1.2300 4.0450 1.3800 ;
        RECT  3.0650 1.2900 3.9050 1.4100 ;
        RECT  3.7450 0.3800 3.8650 1.4100 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5300 0.8700 8.6500 1.3300 ;
        RECT  8.4800 0.8850 8.6500 1.3200 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8000 1.1250 9.0500 1.3100 ;
        RECT  8.7700 0.8850 8.9200 1.2500 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1450 1.2300 10.3500 1.4700 ;
        RECT  9.8700 1.2300 10.3500 1.3800 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5500 0.8700 10.6700 1.1100 ;
        RECT  9.6300 0.9700 10.6700 1.0900 ;
        RECT  10.0100 0.9400 10.4250 1.0900 ;
        RECT  10.0100 0.8700 10.1300 1.1100 ;
        RECT  9.4100 1.2600 9.7500 1.3800 ;
        RECT  9.6300 0.9700 9.7500 1.3800 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5700 0.7400 0.8100 0.8600 ;
        RECT  0.6500 0.7400 0.8000 1.1450 ;
        RECT  0.6500 0.7400 0.7700 1.4200 ;
        RECT  0.6300 1.3000 0.7500 1.9900 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9800 0.6800 2.1000 1.5850 ;
        RECT  1.9200 1.3400 2.0400 1.9900 ;
        RECT  1.8100 1.4650 2.0400 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.4900 -0.1800 10.6100 0.7500 ;
        RECT  8.9900 -0.1800 9.1100 0.7500 ;
        RECT  6.8000 -0.1800 6.9200 0.6300 ;
        RECT  5.3600 0.5900 5.6000 0.7100 ;
        RECT  5.4800 -0.1800 5.6000 0.7100 ;
        RECT  2.9650 -0.1800 3.0850 0.8900 ;
        RECT  1.5000 -0.1800 1.6200 0.7300 ;
        RECT  0.1500 -0.1800 0.2700 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.3100 1.8800 10.4300 2.7900 ;
        RECT  9.0300 1.8800 9.1500 2.7900 ;
        RECT  6.9000 2.1100 7.0200 2.7900 ;
        RECT  5.8800 2.2900 6.1200 2.7900 ;
        RECT  3.6300 2.0300 3.8700 2.1500 ;
        RECT  3.6300 2.0300 3.7500 2.7900 ;
        RECT  2.8500 1.9700 2.9700 2.7900 ;
        RECT  1.5000 1.3400 1.6200 2.7900 ;
        RECT  0.2100 1.3400 0.3300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.0300 0.7500 10.9100 0.7500 10.9100 1.8300 10.8500 1.8300 10.8500 2.0000
                 10.7300 2.0000 10.7300 1.7100 9.8700 1.7100 9.8700 1.6200 9.7500 1.6200 9.7500 1.5000
                 9.9900 1.5000 9.9900 1.5900 10.7900 1.5900 10.7900 0.6300 10.9100 0.6300
                 10.9100 0.5100 11.0300 0.5100 ;
        POLYGON  9.9700 0.7500 9.5100 0.7500 9.5100 0.9900 9.2900 0.9900 9.2900 1.5700 9.6300 1.5700
                 9.6300 1.8300 9.7900 1.8300 9.7900 2.0700 9.6700 2.0700 9.6700 1.9500 9.5100 1.9500
                 9.5100 1.6900 8.1200 1.6900 8.1200 1.5700 8.2400 1.5700 8.2400 0.7200 8.1200 0.7200
                 8.1200 0.6000 8.3600 0.6000 8.3600 1.5700 9.1700 1.5700 9.1700 0.8700 9.3900 0.8700
                 9.3900 0.6300 9.8500 0.6300 9.8500 0.5100 9.9700 0.5100 ;
        POLYGON  8.7900 1.9900 7.6200 1.9900 7.6200 2.1500 7.3800 2.1500 7.3800 1.9900 6.5950 1.9900
                 6.5950 2.1700 5.5600 2.1700 5.5600 2.0500 6.4750 2.0500 6.4750 1.8700 7.8800 1.8700
                 7.8800 0.3600 8.6900 0.3600 8.6900 0.7500 8.5700 0.7500 8.5700 0.4800 8.0000 0.4800
                 8.0000 1.8700 8.7900 1.8700 ;
        POLYGON  7.7600 1.3500 7.7200 1.3500 7.7200 1.7500 7.6000 1.7500 7.6000 1.3500 6.6000 1.3500
                 6.6000 1.2300 7.6400 1.2300 7.6400 0.5400 7.7600 0.5400 ;
        POLYGON  7.5200 1.0600 7.2800 1.0600 7.2800 0.8700 6.5600 0.8700 6.5600 0.5000 6.2000 0.5000
                 6.2000 0.7200 6.0800 0.7200 6.0800 1.1900 5.6400 1.1900 5.6400 1.6900 5.4000 1.6900
                 5.4000 1.5700 5.5200 1.5700 5.5200 1.1900 4.6450 1.1900 4.6450 1.0300 4.8800 1.0300
                 4.8800 0.6200 5.0000 0.6200 5.0000 1.0700 5.9600 1.0700 5.9600 0.6000 6.0800 0.6000
                 6.0800 0.3800 6.6800 0.3800 6.6800 0.7500 7.4000 0.7500 7.4000 0.9400 7.5200 0.9400 ;
        POLYGON  7.1600 1.1100 6.4800 1.1100 6.4800 1.5100 6.5400 1.5100 6.5400 1.7500 6.0100 1.7500
                 6.0100 1.9300 5.0700 1.9300 5.0700 1.4300 4.4050 1.4300 4.4050 0.7100 4.6450 0.7100
                 4.6450 0.8300 4.5250 0.8300 4.5250 1.3100 5.1900 1.3100 5.1900 1.8100 5.8900 1.8100
                 5.8900 1.6300 6.3600 1.6300 6.3600 1.1100 6.3200 1.1100 6.3200 0.6200 6.4400 0.6200
                 6.4400 0.9900 7.1600 0.9900 ;
        POLYGON  4.7700 1.8500 4.6500 1.8500 4.6500 1.6700 2.7100 1.6700 2.7100 1.5500 4.1650 1.5500
                 4.1650 0.8300 3.9850 0.8300 3.9850 0.7100 4.2850 0.7100 4.2850 1.5500 4.7700 1.5500 ;
        POLYGON  4.4100 1.9100 3.4950 1.9100 3.4950 2.0300 3.2100 2.0300 3.2100 1.9100 3.3750 1.9100
                 3.3750 1.7900 4.4100 1.7900 ;
        POLYGON  3.6250 1.1700 2.5900 1.1700 2.5900 1.9100 2.6100 1.9100 2.6100 2.0300 2.3700 2.0300
                 2.3700 1.9100 2.4700 1.9100 2.4700 0.7700 2.5450 0.7700 2.5450 0.6500 2.5350 0.6500
                 2.5350 0.5600 1.8600 0.5600 1.8600 1.1800 1.6200 1.1800 1.6200 1.0600 1.7400 1.0600
                 1.7400 0.4400 2.6550 0.4400 2.6550 0.5300 2.6650 0.5300 2.6650 0.8900 2.5900 0.8900
                 2.5900 1.0500 3.6250 1.0500 ;
        POLYGON  1.1400 1.5800 1.0200 1.5800 1.0200 0.6200 0.4500 0.6200 0.4500 1.0600 0.5300 1.0600
                 0.5300 1.1800 0.2900 1.1800 0.2900 1.0600 0.3300 1.0600 0.3300 0.5000 1.1400 0.5000 ;
    END
END SDFFSX1

MACRO SDFFSRXL
    CLASS CORE ;
    FOREIGN SDFFSRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.7600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 1.5050 2.1750 1.7300 ;
        RECT  1.7550 1.4200 2.0150 1.6700 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9250 2.1100 7.8050 2.2300 ;
        RECT  6.9250 1.8000 7.0450 2.2300 ;
        RECT  5.2950 1.8000 7.0450 1.9200 ;
        RECT  5.2950 1.4400 5.4150 1.9200 ;
        RECT  3.5650 1.4400 5.4150 1.5600 ;
        RECT  3.5650 1.2300 3.7550 1.5600 ;
        RECT  3.4450 1.2600 3.7550 1.3800 ;
        RECT  3.4950 1.2300 3.7550 1.3800 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.0550 1.5200 10.5850 1.6400 ;
        RECT  10.0550 1.5200 10.4750 1.6700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.8050 1.2400 10.9250 1.4800 ;
        RECT  10.4550 1.2400 10.9250 1.3800 ;
        RECT  10.4550 1.2300 10.7150 1.3800 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.8450 1.2200 12.1800 1.4300 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 0.9400 12.4550 1.0900 ;
        RECT  12.3000 0.8700 12.4200 1.1100 ;
        RECT  11.2850 0.9800 12.4200 1.1000 ;
        RECT  11.6050 0.8500 11.7250 1.1000 ;
        RECT  11.2850 0.9800 11.4050 1.6700 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1500 1.3400 0.2700 1.5800 ;
        RECT  0.1350 0.6800 0.2550 0.9600 ;
        RECT  0.1300 0.8400 0.2500 1.4600 ;
        RECT  0.0700 0.8850 0.2500 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4150 1.5850 1.5350 2.0900 ;
        RECT  1.4150 0.6800 1.5350 0.9600 ;
        RECT  1.2300 1.4650 1.4950 1.7250 ;
        RECT  1.3750 0.8400 1.4950 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.7600 0.1800 ;
        RECT  12.0850 -0.1800 12.2050 0.7500 ;
        RECT  10.6850 0.5000 10.9250 0.6200 ;
        RECT  10.8050 -0.1800 10.9250 0.6200 ;
        RECT  9.6950 -0.1800 9.9350 0.3200 ;
        RECT  7.8250 -0.1800 7.9450 0.8600 ;
        RECT  3.1250 -0.1800 3.3650 0.3200 ;
        RECT  1.8350 -0.1800 1.9550 0.9200 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.7600 2.7900 ;
        RECT  12.0850 1.9700 12.2050 2.7900 ;
        RECT  10.7450 2.0300 10.9850 2.1500 ;
        RECT  10.7450 2.0300 10.8650 2.7900 ;
        RECT  9.8750 2.0300 10.1150 2.1500 ;
        RECT  9.8750 2.0300 9.9950 2.7900 ;
        RECT  7.9450 2.2300 8.0650 2.7900 ;
        RECT  6.2250 2.2900 6.4650 2.7900 ;
        RECT  4.4450 2.1600 4.6850 2.2800 ;
        RECT  4.4450 2.1600 4.5650 2.7900 ;
        RECT  3.1850 2.1700 3.3050 2.7900 ;
        RECT  1.8350 1.9700 1.9550 2.7900 ;
        RECT  0.5700 1.4600 0.6900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.6950 1.7900 12.6250 1.7900 12.6250 2.0900 12.5050 2.0900 12.5050 1.6700
                 11.6050 1.6700 11.6050 1.4300 11.7250 1.4300 11.7250 1.5500 12.5750 1.5500
                 12.5750 0.6900 12.4450 0.6900 12.4450 0.5700 12.6950 0.5700 ;
        POLYGON  11.6250 0.6900 11.4300 0.6900 11.4300 0.8600 11.1650 0.8600 11.1650 1.7900
                 11.5650 1.7900 11.5650 2.0900 11.4450 2.0900 11.4450 1.9100 11.0450 1.9100
                 11.0450 0.8600 10.4450 0.8600 10.4450 0.5600 9.0050 0.5600 9.0050 0.7400 9.0650 0.7400
                 9.0650 1.5800 9.1850 1.5800 9.1850 1.8200 9.0650 1.8200 9.0650 1.7000 8.9450 1.7000
                 8.9450 0.8600 8.8850 0.8600 8.8850 0.4400 10.5650 0.4400 10.5650 0.7400 11.3100 0.7400
                 11.3100 0.5700 11.6250 0.5700 ;
        POLYGON  10.5050 2.0900 10.3850 2.0900 10.3850 1.9100 9.6700 1.9100 9.6700 2.0600 8.6850 2.0600
                 8.6850 2.2000 8.4450 2.2000 8.4450 2.0600 7.9600 2.0600 7.9600 1.9900 7.1650 1.9900
                 7.1650 1.6000 6.7350 1.6000 6.7350 1.4100 6.6150 1.4100 6.6150 1.2900 6.8550 1.2900
                 6.8550 1.4800 7.2850 1.4800 7.2850 1.8700 8.0800 1.8700 8.0800 1.9400 9.5500 1.9400
                 9.5500 1.7900 9.8150 1.7900 9.8150 1.1100 9.6650 1.1100 9.6650 1.2000 9.5450 1.2000
                 9.5450 0.9600 9.6650 0.9600 9.6650 0.9900 10.0850 0.9900 10.0850 0.6800 10.3250 0.6800
                 10.3250 0.8000 10.2050 0.8000 10.2050 1.1100 9.9350 1.1100 9.9350 1.7900
                 10.5050 1.7900 ;
        POLYGON  9.6350 1.6700 9.3050 1.6700 9.3050 1.4000 9.1850 1.4000 9.1850 1.1600 9.2150 1.1600
                 9.2150 0.6800 9.4550 0.6800 9.4550 0.8000 9.3350 0.8000 9.3350 1.2800 9.4250 1.2800
                 9.4250 1.5500 9.6350 1.5500 ;
        POLYGON  8.8250 1.7600 8.5850 1.7600 8.5850 1.1200 7.2650 1.1200 7.2650 1.0000 8.4650 1.0000
                 8.4650 0.6200 8.5850 0.6200 8.5850 1.0000 8.7050 1.0000 8.7050 1.6400 8.8250 1.6400 ;
        POLYGON  8.1450 1.3600 7.5250 1.3600 7.5250 1.6300 7.6450 1.6300 7.6450 1.7500 7.4050 1.7500
                 7.4050 1.3600 6.9850 1.3600 6.9850 1.0400 6.4950 1.0400 6.4950 1.6800 5.9550 1.6800
                 5.9550 1.5600 6.3750 1.5600 6.3750 1.0400 6.0550 1.0400 6.0550 0.6600 6.1750 0.6600
                 6.1750 0.9200 6.9850 0.9200 6.9850 0.6200 7.1050 0.6200 7.1050 1.2400 8.1450 1.2400 ;
        POLYGON  7.5250 0.8600 7.4050 0.8600 7.4050 0.6200 7.2250 0.6200 7.2250 0.5000 6.7450 0.5000
                 6.7450 0.8000 6.5050 0.8000 6.5050 0.6800 6.6250 0.6800 6.6250 0.3800 7.3450 0.3800
                 7.3450 0.5000 7.5250 0.5000 ;
        POLYGON  6.8050 2.1700 6.5500 2.1700 6.5500 2.1600 4.9600 2.1600 4.9600 2.0400 4.2850 2.0400
                 4.2850 2.2500 4.1650 2.2500 4.1650 2.0400 3.1700 2.0400 3.1700 2.0500 2.3750 2.0500
                 2.3750 2.0900 2.2550 2.0900 2.2550 1.8500 2.3150 1.8500 2.3150 0.6800 2.4350 0.6800
                 2.4350 1.9300 3.0500 1.9300 3.0500 1.9200 5.0800 1.9200 5.0800 2.0400 6.6700 2.0400
                 6.6700 2.0500 6.8050 2.0500 ;
        POLYGON  6.2550 1.3600 5.8150 1.3600 5.8150 0.5200 5.3750 0.5200 5.3750 0.4000 5.9350 0.4000
                 5.9350 1.2400 6.2550 1.2400 ;
        POLYGON  5.7750 1.6800 5.5350 1.6800 5.5350 1.5600 5.5750 1.5600 5.5750 1.3200 4.2250 1.3200
                 4.2250 1.1100 3.3250 1.1100 3.3250 1.1800 2.9050 1.1800 2.9050 1.0600 3.2050 1.0600
                 3.2050 0.9900 4.3450 0.9900 4.3450 1.2000 5.5750 1.2000 5.5750 0.6600 5.6950 0.6600
                 5.6950 1.5600 5.7750 1.5600 ;
        POLYGON  5.2750 0.9000 5.1850 0.9000 5.1850 1.0800 4.4650 1.0800 4.4650 0.8400 4.2850 0.8400
                 4.2850 0.7200 4.5850 0.7200 4.5850 0.9600 5.0650 0.9600 5.0650 0.7800 5.1550 0.7800
                 5.1550 0.6600 5.2750 0.6600 ;
        RECT  3.6050 1.6800 5.1750 1.8000 ;
        POLYGON  4.9450 0.8400 4.7050 0.8400 4.7050 0.6000 4.1650 0.6000 4.1650 0.7600 3.8450 0.7600
                 3.8450 0.8400 3.6050 0.8400 3.6050 0.7200 3.7250 0.7200 3.7250 0.6400 4.0450 0.6400
                 4.0450 0.4800 4.8250 0.4800 4.8250 0.7200 4.9450 0.7200 ;
        POLYGON  3.9250 0.5200 3.6050 0.5200 3.6050 0.5600 2.8250 0.5600 2.8250 0.9000 2.7850 0.9000
                 2.7850 1.5700 2.8250 1.5700 2.8250 1.8100 2.7050 1.8100 2.7050 1.6900 2.6650 1.6900
                 2.6650 0.7800 2.7050 0.7800 2.7050 0.5600 2.1950 0.5600 2.1950 1.2000 1.6150 1.2000
                 1.6150 1.0800 2.0750 1.0800 2.0750 0.4400 3.4850 0.4400 3.4850 0.4000 3.9250 0.4000 ;
        POLYGON  1.1450 1.0800 1.1100 1.0800 1.1100 1.5800 0.9900 1.5800 0.9900 1.2000 0.3700 1.2000
                 0.3700 1.0800 0.9900 1.0800 0.9900 0.9600 1.0250 0.9600 1.0250 0.6800 1.1450 0.6800 ;
    END
END SDFFSRXL

MACRO SDFFSRX4
    CLASS CORE ;
    FOREIGN SDFFSRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 16.5300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6550 1.4600 1.8950 1.5800 ;
        RECT  1.6550 0.3600 1.7750 1.5800 ;
        RECT  0.9550 0.3600 1.7750 0.4800 ;
        RECT  0.3550 0.9200 1.2950 1.0400 ;
        RECT  0.8850 0.9200 1.1450 1.0900 ;
        RECT  0.9550 0.3600 1.0750 1.0900 ;
        RECT  0.3550 0.9200 0.4750 1.1600 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2350 0.9550 1.4350 ;
        RECT  0.5950 1.2100 0.8550 1.4350 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.9350 1.1750 2.2500 1.2950 ;
        RECT  1.9350 1.0550 2.0550 1.2950 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9000 2.8850 1.1200 ;
        RECT  2.6550 0.9000 2.7750 1.2900 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9750 1.1650 7.2350 1.3800 ;
        RECT  7.1050 1.0000 7.2250 1.3800 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5550 1.1850 7.8150 1.3800 ;
        RECT  7.5650 1.0000 7.6850 1.3800 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1650 0.7000 13.3650 0.8200 ;
        RECT  13.1850 1.4400 13.3050 2.2100 ;
        RECT  12.9050 1.4400 13.3050 1.5600 ;
        RECT  12.2500 1.3200 13.0250 1.4400 ;
        RECT  12.2800 0.7000 12.4000 1.5600 ;
        RECT  12.2450 1.4400 12.3650 2.2100 ;
        RECT  12.2500 1.1750 12.4000 1.5600 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  14.0850 0.7000 15.2850 0.8200 ;
        RECT  14.9050 1.5600 15.0250 2.2100 ;
        RECT  14.8850 1.3200 15.0050 1.6800 ;
        RECT  14.2450 1.3200 15.0050 1.4400 ;
        RECT  14.2450 1.1750 14.4300 1.4400 ;
        RECT  14.0650 1.4400 14.3650 1.5600 ;
        RECT  14.2450 0.7000 14.3650 1.5600 ;
        RECT  14.0650 1.4400 14.1850 2.2100 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 16.5300 0.1800 ;
        RECT  15.6450 0.5100 15.8850 0.6300 ;
        RECT  15.7650 -0.1800 15.8850 0.6300 ;
        RECT  14.5650 -0.1800 14.8050 0.3400 ;
        RECT  13.6050 -0.1800 13.8450 0.3400 ;
        RECT  12.6450 -0.1800 12.8850 0.3400 ;
        RECT  11.5650 0.6000 11.8050 0.7200 ;
        RECT  11.5650 -0.1800 11.6850 0.7200 ;
        RECT  10.7850 -0.1800 10.9050 0.8600 ;
        RECT  7.3050 0.5200 7.5450 0.6400 ;
        RECT  7.3050 -0.1800 7.4250 0.6400 ;
        RECT  4.7050 -0.1800 4.9450 0.3400 ;
        RECT  1.8950 -0.1800 2.0150 0.7800 ;
        RECT  0.6150 -0.1800 0.7350 0.7800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 16.5300 2.7900 ;
        RECT  15.3250 1.5600 15.4450 2.7900 ;
        RECT  14.4850 1.5600 14.6050 2.7900 ;
        RECT  13.6450 1.5600 13.7650 2.7900 ;
        RECT  12.6650 1.5600 12.7850 2.7900 ;
        RECT  11.8250 1.6000 11.9450 2.7900 ;
        RECT  10.9850 1.7600 11.1050 2.7900 ;
        RECT  9.9250 1.8800 10.0450 2.7900 ;
        RECT  7.2150 1.9800 7.3350 2.7900 ;
        RECT  7.0950 1.9800 7.3350 2.1000 ;
        RECT  5.4350 2.2400 5.6750 2.7900 ;
        RECT  4.5650 2.2400 4.8050 2.7900 ;
        RECT  2.1550 1.9400 2.3950 2.0600 ;
        RECT  2.1550 1.9400 2.2750 2.7900 ;
        RECT  0.6750 1.8800 0.7950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  16.2450 1.4400 15.8650 1.4400 15.8650 2.2100 15.7450 2.2100 15.7450 1.4400
                 15.1250 1.4400 15.1250 1.3000 15.3650 1.3000 15.3650 1.3200 16.1250 1.3200
                 16.1250 0.6400 16.2450 0.6400 ;
        POLYGON  15.7250 1.2000 15.6050 1.2000 15.6050 0.8700 15.4050 0.8700 15.4050 0.5800
                 12.0450 0.5800 12.0450 0.9600 11.5050 0.9600 11.5050 1.2200 12.1250 1.2200
                 12.1250 1.3400 11.5250 1.3400 11.5250 2.1200 11.4050 2.1200 11.4050 1.3400
                 11.3850 1.3400 11.3850 1.1400 10.2450 1.1400 10.2450 1.0200 11.2050 1.0200
                 11.2050 0.6400 11.3250 0.6400 11.3250 0.8400 11.9250 0.8400 11.9250 0.4600
                 15.5250 0.4600 15.5250 0.7500 15.7250 0.7500 ;
        POLYGON  11.2650 1.5200 8.8450 1.5200 8.8450 1.8900 8.7250 1.8900 8.7250 1.4000 8.6550 1.4000
                 8.6550 0.6800 8.7750 0.6800 8.7750 1.2800 8.8450 1.2800 8.8450 1.4000 11.1450 1.4000
                 11.1450 1.2600 11.2650 1.2600 ;
        POLYGON  10.7450 1.9400 10.2650 1.9400 10.2650 1.7600 9.5900 1.7600 9.5900 1.8100 9.0850 1.8100
                 9.0850 1.6900 9.4700 1.6900 9.4700 1.6400 10.3850 1.6400 10.3850 1.8200 10.7450 1.8200 ;
        POLYGON  10.4850 0.8600 10.3650 0.8600 10.3650 0.7400 10.1850 0.7400 10.1850 0.5000
                 9.7750 0.5000 9.7750 0.8000 9.4650 0.8000 9.4650 0.6800 9.6550 0.6800 9.6550 0.3800
                 10.3050 0.3800 10.3050 0.6200 10.4850 0.6200 ;
        POLYGON  10.0650 1.0400 9.2250 1.0400 9.2250 0.9200 9.1350 0.9200 9.1350 0.6800 9.2550 0.6800
                 9.2550 0.8000 9.3450 0.8000 9.3450 0.9200 9.9450 0.9200 9.9450 0.6200 10.0650 0.6200 ;
        POLYGON  9.8650 1.2800 8.9850 1.2800 8.9850 1.1600 8.8950 1.1600 8.8950 0.5600 7.9650 0.5600
                 7.9650 0.7400 8.0550 0.7400 8.0550 1.6200 7.9350 1.6200 7.9350 0.8600 7.7850 0.8600
                 7.7850 0.8800 7.0650 0.8800 7.0650 0.5000 6.6500 0.5000 6.6500 0.4800 6.2650 0.4800
                 6.2650 0.3600 6.7700 0.3600 6.7700 0.3800 7.1850 0.3800 7.1850 0.7600 7.6650 0.7600
                 7.6650 0.6200 7.8450 0.6200 7.8450 0.4400 9.0150 0.4400 9.0150 1.0400 9.1050 1.0400
                 9.1050 1.1600 9.8650 1.1600 ;
        POLYGON  9.1050 2.2500 7.9550 2.2500 7.9550 2.1300 7.4550 2.1300 7.4550 1.8600 6.3750 1.8600
                 6.3750 1.6400 5.0450 1.6400 5.0450 1.5200 5.1850 1.5200 5.1850 1.0000 4.3450 1.0000
                 4.3450 1.2800 4.2250 1.2800 4.2250 0.8800 5.1850 0.8800 5.1850 0.7000 5.4250 0.7000
                 5.4250 0.8200 5.3050 0.8200 5.3050 1.5200 6.4950 1.5200 6.4950 1.7400 7.5750 1.7400
                 7.5750 2.0100 8.0750 2.0100 8.0750 2.1300 8.4850 2.1300 8.4850 1.6400 8.4150 1.6400
                 8.4150 1.0400 8.5350 1.0400 8.5350 1.5200 8.6050 1.5200 8.6050 2.1300 9.1050 2.1300 ;
        POLYGON  8.3650 2.0100 8.2450 2.0100 8.2450 1.8900 7.6950 1.8900 7.6950 1.6200 6.6150 1.6200
                 6.6150 1.4000 5.5450 1.4000 5.5450 0.5800 4.4650 0.5800 4.4650 0.5000 4.3450 0.5000
                 4.3450 0.3800 4.5850 0.3800 4.5850 0.4600 5.5250 0.4600 5.5250 0.3800 6.1450 0.3800
                 6.1450 0.6000 6.4650 0.6000 6.4650 0.6800 6.5850 0.6800 6.5850 0.8000 6.3450 0.8000
                 6.3450 0.7200 6.0250 0.7200 6.0250 0.5000 5.6650 0.5000 5.6650 1.2800 6.8550 1.2800
                 6.8550 1.5000 7.8150 1.5000 7.8150 1.7700 8.1750 1.7700 8.1750 0.8000 8.2350 0.8000
                 8.2350 0.6800 8.3550 0.6800 8.3550 0.9200 8.2950 0.9200 8.2950 1.7700 8.3650 1.7700 ;
        POLYGON  6.9750 2.2500 6.4000 2.2500 6.4000 2.1000 6.1350 2.1000 6.1350 1.8800 4.8050 1.8800
                 4.8050 1.5200 4.2450 1.5200 4.2450 1.5600 4.0050 1.5600 4.0050 1.5200 3.9850 1.5200
                 3.9850 0.5200 3.5000 0.5200 3.5000 0.5400 2.5550 0.5400 2.5550 0.6600 3.1250 0.6600
                 3.1250 1.9400 2.7550 1.9400 2.7550 1.8200 3.0050 1.8200 3.0050 0.7800 2.4350 0.7800
                 2.4350 0.4200 3.3800 0.4200 3.3800 0.4000 3.5250 0.4000 3.5250 0.3600 3.7650 0.3600
                 3.7650 0.4000 4.1050 0.4000 4.1050 1.4000 4.8050 1.4000 4.8050 1.1200 4.9650 1.1200
                 4.9650 1.3600 4.9250 1.3600 4.9250 1.7600 6.2550 1.7600 6.2550 1.9800 6.5200 1.9800
                 6.5200 2.1300 6.9750 2.1300 ;
        POLYGON  6.9450 1.0400 5.7850 1.0400 5.7850 0.6200 5.9050 0.6200 5.9050 0.9200 6.8250 0.9200
                 6.8250 0.6200 6.9450 0.6200 ;
        POLYGON  6.0150 2.1200 4.4500 2.1200 4.4500 2.0600 3.9250 2.0600 3.9250 1.8200 3.7450 1.8200
                 3.7450 0.6400 3.8650 0.6400 3.8650 1.7000 4.0450 1.7000 4.0450 1.9400 4.5700 1.9400
                 4.5700 2.0000 6.0150 2.0000 ;
        POLYGON  3.6250 2.1800 2.5150 2.1800 2.5150 1.8200 1.5750 1.8200 1.5750 2.0000 1.4550 2.0000
                 1.4550 1.8800 1.4150 1.8800 1.4150 0.7200 1.1950 0.7200 1.1950 0.6000 1.5350 0.6000
                 1.5350 1.7000 2.6350 1.7000 2.6350 2.0600 3.5050 2.0600 3.5050 0.8200 3.2650 0.8200
                 3.2650 0.7000 3.6250 0.7000 ;
        POLYGON  1.2950 1.6750 0.3750 1.6750 0.3750 2.0000 0.2550 2.0000 0.2550 1.7950 0.1150 1.7950
                 0.1150 0.6800 0.1950 0.6800 0.1950 0.5400 0.3150 0.5400 0.3150 0.8000 0.2350 0.8000
                 0.2350 1.5550 1.1750 1.5550 1.1750 1.2100 1.2950 1.2100 ;
    END
END SDFFSRX4

MACRO SDFFSRX2
    CLASS CORE ;
    FOREIGN SDFFSRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 15.0800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5750 0.3600 1.6950 1.7000 ;
        RECT  0.8950 0.3600 1.6950 0.4800 ;
        RECT  0.9750 0.9400 1.2150 1.0600 ;
        RECT  0.3900 0.9000 1.0950 1.0200 ;
        RECT  0.8950 0.3600 1.0150 1.0200 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        RECT  0.3900 0.9000 0.5100 1.4350 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 1.1400 0.8550 1.5700 ;
        RECT  0.6500 1.1400 0.8550 1.5550 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 0.8850 2.2500 1.1450 ;
        RECT  1.8150 0.9000 2.2500 1.0200 ;
        RECT  1.8150 0.9000 1.9350 1.1400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0350 2.5400 1.5000 ;
        RECT  2.3900 0.9600 2.5100 1.5000 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.8760  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 7.3000  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 0.9450 5.3300 1.1200 ;
        RECT  4.9450 0.9400 5.2050 1.1400 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 1.1200 12.4550 1.3800 ;
        RECT  12.1850 1.1000 12.4250 1.3400 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.9050 0.6800 13.0250 2.0300 ;
        RECT  12.8300 1.4650 13.0250 1.7250 ;
        RECT  12.8600 1.3800 13.0250 1.7250 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.7250 0.7400 14.0450 0.8600 ;
        RECT  13.7450 1.3000 13.8650 2.0300 ;
        RECT  13.7250 0.7400 13.8450 1.4200 ;
        RECT  13.4100 1.0250 13.8450 1.1450 ;
        RECT  13.4100 0.8850 13.5600 1.1450 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 15.0800 0.1800 ;
        RECT  14.2850 -0.1800 14.5250 0.3200 ;
        RECT  13.3250 -0.1800 13.5650 0.3200 ;
        RECT  12.3650 -0.1800 12.6050 0.3200 ;
        RECT  11.2100 -0.1800 11.3300 0.8300 ;
        RECT  4.9900 -0.1800 5.2300 0.3200 ;
        RECT  2.9000 -0.1800 3.0200 0.9200 ;
        RECT  1.8600 -0.1800 1.9800 0.7800 ;
        RECT  0.5550 -0.1800 0.6750 0.7800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 15.0800 2.7900 ;
        RECT  14.1650 1.3800 14.2850 2.7900 ;
        RECT  13.3250 1.3800 13.4450 2.7900 ;
        RECT  12.4850 1.5000 12.6050 2.7900 ;
        RECT  10.9500 2.1300 11.0700 2.7900 ;
        RECT  10.8300 2.1300 11.0700 2.2500 ;
        RECT  8.4500 1.8800 8.5700 2.7900 ;
        RECT  8.3300 1.8800 8.5700 2.0000 ;
        RECT  6.2300 1.9600 6.3500 2.7900 ;
        RECT  6.1100 1.9600 6.3500 2.0800 ;
        RECT  4.8500 2.1300 4.9700 2.7900 ;
        RECT  2.9250 2.2800 3.1650 2.7900 ;
        RECT  2.0550 1.8600 2.1750 2.7900 ;
        RECT  0.6950 1.9300 0.8150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  15.0050 0.8600 14.8850 0.8600 14.8850 1.1800 14.7050 1.1800 14.7050 1.6200
                 14.5850 1.6200 14.5850 1.1800 13.9650 1.1800 13.9650 1.0600 14.7650 1.0600
                 14.7650 0.7400 15.0050 0.7400 ;
        POLYGON  14.8850 0.5200 14.7650 0.5200 14.7650 0.5600 13.2650 0.5600 13.2650 1.2600
                 13.1450 1.2600 13.1450 0.5600 12.7850 0.5600 12.7850 1.2600 12.6650 1.2600
                 12.6650 0.6000 11.7500 0.6000 11.7500 0.8400 11.7100 0.8400 11.7100 1.5900
                 11.5500 1.5900 11.5500 2.0100 11.4300 2.0100 11.4300 1.4700 11.5900 1.4700
                 11.5900 1.1100 10.4900 1.1100 10.4900 0.9900 11.5900 0.9900 11.5900 0.7200
                 11.6300 0.7200 11.6300 0.4800 12.6650 0.4800 12.6650 0.4400 14.6450 0.4400
                 14.6450 0.4000 14.8850 0.4000 ;
        POLYGON  12.2000 0.8400 12.0650 0.8400 12.0650 1.6200 12.1850 1.6200 12.1850 2.2500
                 11.1900 2.2500 11.1900 2.0100 8.9300 2.0100 8.9300 1.5200 8.1100 1.5200 8.1100 1.4000
                 9.0500 1.4000 9.0500 1.8900 11.3100 1.8900 11.3100 2.1300 12.0650 2.1300
                 12.0650 1.7400 11.9450 1.7400 11.9450 0.7200 12.2000 0.7200 ;
        POLYGON  11.4700 1.3500 9.4100 1.3500 9.4100 1.0400 7.6100 1.0400 7.6100 1.6000 7.5500 1.6000
                 7.5500 1.7200 7.4300 1.7200 7.4300 1.4800 7.4900 1.4800 7.4900 0.6200 7.6100 0.6200
                 7.6100 0.9200 9.5300 0.9200 9.5300 1.2300 11.4700 1.2300 ;
        POLYGON  10.9100 0.8300 10.7900 0.8300 10.7900 0.5900 10.6700 0.5900 10.6700 0.5300
                 10.1300 0.5300 10.1300 0.7700 9.8900 0.7700 9.8900 0.6500 10.0100 0.6500
                 10.0100 0.4100 10.7900 0.4100 10.7900 0.4700 10.9100 0.4700 ;
        POLYGON  10.7100 2.2500 8.6900 2.2500 8.6900 1.7600 8.2100 1.7600 8.2100 1.9600 7.6800 1.9600
                 7.6800 2.2000 6.4700 2.2000 6.4700 1.8400 5.9900 1.8400 5.9900 2.2500 5.1100 2.2500
                 5.1100 2.1300 5.8700 2.1300 5.8700 1.7200 6.5900 1.7200 6.5900 2.0800 7.5600 2.0800
                 7.5600 1.8400 8.0900 1.8400 8.0900 1.6400 8.8100 1.6400 8.8100 2.1300 10.7100 2.1300 ;
        POLYGON  10.5900 1.7700 9.1700 1.7700 9.1700 1.2800 7.9900 1.2800 7.9900 1.5200 7.9700 1.5200
                 7.9700 1.7200 7.8500 1.7200 7.8500 1.4000 7.8700 1.4000 7.8700 1.1600 9.2900 1.1600
                 9.2900 1.6500 10.5900 1.6500 ;
        POLYGON  10.5500 0.7700 10.3700 0.7700 10.3700 1.0100 9.6500 1.0100 9.6500 0.8000 7.8500 0.8000
                 7.8500 0.6800 9.7700 0.6800 9.7700 0.8900 10.2500 0.8900 10.2500 0.6500 10.5500 0.6500 ;
        POLYGON  7.8100 0.4800 7.3700 0.4800 7.3700 1.2800 7.3100 1.2800 7.3100 1.9600 6.7100 1.9600
                 6.7100 1.6000 5.7500 1.6000 5.7500 2.0100 4.9600 2.0100 4.9600 1.6200 4.4300 1.6200
                 4.4300 1.1400 4.5500 1.1400 4.5500 1.5000 5.0800 1.5000 5.0800 1.8900 5.6300 1.8900
                 5.6300 1.4800 6.8300 1.4800 6.8300 1.8400 7.1900 1.8400 7.1900 1.1600 7.2500 1.1600
                 7.2500 0.3600 7.8100 0.3600 ;
        POLYGON  7.1300 1.0400 7.0700 1.0400 7.0700 1.7200 6.9500 1.7200 6.9500 1.3600 5.4450 1.3600
                 5.4450 1.6500 5.5100 1.6500 5.5100 1.7700 5.2700 1.7700 5.2700 1.6500 5.3250 1.6500
                 5.3250 1.3800 4.7300 1.3800 4.7300 1.2600 5.3250 1.2600 5.3250 1.2400 6.1700 1.2400
                 6.1700 0.6200 6.2900 0.6200 6.2900 1.2400 6.9500 1.2400 6.9500 0.9200 7.0100 0.9200
                 7.0100 0.6200 7.1300 0.6200 ;
        POLYGON  6.7100 0.8600 6.5900 0.8600 6.5900 0.7400 6.4600 0.7400 6.4600 0.5000 6.0500 0.5000
                 6.0500 0.8000 5.6900 0.8000 5.6900 0.6800 5.9300 0.6800 5.9300 0.3800 6.5800 0.3800
                 6.5800 0.6200 6.7100 0.6200 ;
        POLYGON  5.8100 0.4800 5.6900 0.4800 5.6900 0.5600 4.7500 0.5600 4.7500 0.5000 4.0700 0.5000
                 4.0700 1.6300 4.0300 1.6300 4.0300 1.7500 3.9100 1.7500 3.9100 1.5100 3.9500 1.5100
                 3.9500 0.5000 3.4400 0.5000 3.4400 0.8000 3.5500 0.8000 3.5500 1.7000 3.5400 1.7000
                 3.5400 1.8200 3.4200 1.8200 3.4200 1.5800 3.4300 1.5800 3.4300 0.9200 3.3200 0.9200
                 3.3200 0.3800 4.3650 0.3800 4.3650 0.3600 4.6050 0.3600 4.6050 0.3800 4.8700 0.3800
                 4.8700 0.4400 5.5700 0.4400 5.5700 0.3600 5.8100 0.3600 ;
        POLYGON  5.7900 1.1200 5.4500 1.1200 5.4500 0.8200 4.3100 0.8200 4.3100 1.9700 4.2700 1.9700
                 4.2700 2.0900 4.1500 2.0900 4.1500 1.8500 4.1900 1.8500 4.1900 0.6800 4.4300 0.6800
                 4.4300 0.7000 5.5700 0.7000 5.5700 1.0000 5.7900 1.0000 ;
        POLYGON  3.8500 2.2100 3.7300 2.2100 3.7300 2.1600 2.2950 2.1600 2.2950 1.7400 1.9350 1.7400
                 1.9350 1.9400 1.4550 1.9400 1.4550 2.0500 1.3350 2.0500 1.3350 0.7200 1.1350 0.7200
                 1.1350 0.6000 1.4550 0.6000 1.4550 1.8200 1.8150 1.8200 1.8150 1.6200 2.4150 1.6200
                 2.4150 2.0400 3.6700 2.0400 3.6700 0.7400 3.7100 0.7400 3.7100 0.6200 3.8300 0.6200
                 3.8300 0.8600 3.7900 0.8600 3.7900 1.9700 3.8500 1.9700 ;
        POLYGON  3.3100 1.4200 2.7800 1.4200 2.7800 1.9200 2.5350 1.9200 2.5350 1.8000 2.6600 1.8000
                 2.6600 0.7200 2.2550 0.7200 2.2550 0.6000 2.7800 0.6000 2.7800 1.3000 3.3100 1.3000 ;
        POLYGON  1.1950 1.8100 0.3750 1.8100 0.3750 2.0500 0.2550 2.0500 0.2550 1.9300 0.1200 1.9300
                 0.1200 0.9350 0.1350 0.9350 0.1350 0.5400 0.2550 0.5400 0.2550 1.0550 0.2400 1.0550
                 0.2400 1.6900 1.0750 1.6900 1.0750 1.2200 1.1950 1.2200 ;
    END
END SDFFSRX2

MACRO SDFFSRX1
    CLASS CORE ;
    FOREIGN SDFFSRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.7600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.2700 2.2500 1.7250 ;
        RECT  2.1050 1.2500 2.2250 1.7250 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8850 2.1100 7.7650 2.2300 ;
        RECT  6.8850 1.7900 7.0050 2.2300 ;
        RECT  5.2450 1.7900 7.0050 1.9100 ;
        RECT  5.2450 1.4000 5.3650 1.9100 ;
        RECT  3.5150 1.4000 5.3650 1.5200 ;
        RECT  3.5150 1.2300 3.7550 1.5200 ;
        RECT  3.3950 1.2600 3.7550 1.3800 ;
        RECT  3.4950 1.2300 3.7550 1.3800 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.0150 1.5000 10.3650 1.6300 ;
        RECT  9.8750 1.5050 10.1350 1.6700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1650 1.2600 10.7050 1.3800 ;
        RECT  10.1650 1.2300 10.4250 1.3800 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.5850 1.2700 12.0450 1.3900 ;
        RECT  11.6100 1.2300 12.0450 1.3900 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1650 0.9900 12.2850 1.2300 ;
        RECT  11.9050 0.9400 12.1650 1.1100 ;
        RECT  11.0650 0.9900 12.2850 1.1100 ;
        RECT  11.6050 0.8700 11.7250 1.1100 ;
        RECT  11.0650 0.9900 11.1850 1.6300 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4250 1.3200 1.5450 2.0850 ;
        RECT  1.3650 0.6500 1.4850 0.8900 ;
        RECT  1.3250 0.7700 1.4450 1.4400 ;
        RECT  1.2300 0.8850 1.4450 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.7600 0.1800 ;
        RECT  12.0850 -0.1800 12.2050 0.7500 ;
        RECT  10.6850 0.5100 10.9250 0.6300 ;
        RECT  10.8050 -0.1800 10.9250 0.6300 ;
        RECT  9.6950 -0.1800 9.9350 0.3200 ;
        RECT  7.8250 -0.1800 7.9450 0.8600 ;
        RECT  3.0750 -0.1800 3.3150 0.3200 ;
        RECT  1.7850 -0.1800 1.9050 0.8900 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.7600 2.7900 ;
        RECT  11.9050 1.9300 12.0250 2.7900 ;
        RECT  10.5250 1.9900 10.7650 2.1100 ;
        RECT  10.5250 1.9900 10.6450 2.7900 ;
        RECT  9.7150 2.2900 9.9550 2.7900 ;
        RECT  7.9050 2.2300 8.0250 2.7900 ;
        RECT  6.1850 2.2900 6.4250 2.7900 ;
        RECT  4.3950 2.1200 4.6350 2.2400 ;
        RECT  4.3950 2.1200 4.5150 2.7900 ;
        RECT  3.1350 2.1200 3.2550 2.7900 ;
        RECT  1.8450 1.7250 1.9650 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.6850 0.6900 12.5250 0.6900 12.5250 1.7500 12.4450 1.7500 12.4450 2.0500
                 12.3250 2.0500 12.3250 1.6300 11.3450 1.6300 11.3450 1.5100 12.4050 1.5100
                 12.4050 0.5700 12.6850 0.5700 ;
        POLYGON  11.5650 0.7500 11.4850 0.7500 11.4850 0.8700 10.9450 0.8700 10.9450 1.7500
                 11.3450 1.7500 11.3450 2.0500 11.2250 2.0500 11.2250 1.8700 10.8250 1.8700
                 10.8250 0.8700 10.4450 0.8700 10.4450 0.5600 9.0050 0.5600 9.0050 0.7400 9.0250 0.7400
                 9.0250 1.8200 8.9050 1.8200 8.9050 0.8600 8.8850 0.8600 8.8850 0.4400 10.5650 0.4400
                 10.5650 0.7500 11.3650 0.7500 11.3650 0.6300 11.4450 0.6300 11.4450 0.5100
                 11.5650 0.5100 ;
        POLYGON  10.3250 0.8000 10.0450 0.8000 10.0450 1.2000 9.7550 1.2000 9.7550 2.0500
                 10.1650 2.0500 10.1650 1.8400 10.2850 1.8400 10.2850 2.1700 8.5250 2.1700
                 8.5250 2.2000 8.2850 2.2000 8.2850 2.0000 7.8850 2.0000 7.8850 1.9900 7.1250 1.9900
                 7.1250 1.6700 6.7450 1.6700 6.7450 1.4100 6.5650 1.4100 6.5650 1.2900 6.8650 1.2900
                 6.8650 1.5500 7.2450 1.5500 7.2450 1.8700 8.0050 1.8700 8.0050 1.8800 8.4300 1.8800
                 8.4300 2.0500 9.6350 2.0500 9.6350 1.2000 9.5350 1.2000 9.5350 0.9600 9.6550 0.9600
                 9.6550 1.0800 9.9250 1.0800 9.9250 0.6800 10.3250 0.6800 ;
        POLYGON  9.4750 1.9300 9.2350 1.9300 9.2350 1.5000 9.1450 1.5000 9.1450 1.2600 9.2350 1.2600
                 9.2350 0.8000 9.2150 0.8000 9.2150 0.6800 9.4550 0.6800 9.4550 0.8000 9.3550 0.8000
                 9.3550 1.8100 9.4750 1.8100 ;
        POLYGON  8.6650 1.7600 8.4250 1.7600 8.4250 1.6400 8.4650 1.6400 8.4650 1.1900 7.2250 1.1900
                 7.2250 1.0700 8.4650 1.0700 8.4650 0.6200 8.5850 0.6200 8.5850 1.6400 8.6650 1.6400 ;
        POLYGON  8.1450 1.4300 7.4850 1.4300 7.4850 1.6300 7.6050 1.6300 7.6050 1.7500 7.3650 1.7500
                 7.3650 1.4300 6.9850 1.4300 6.9850 1.1700 6.4450 1.1700 6.4450 1.6400 5.9050 1.6400
                 5.9050 1.5200 6.3250 1.5200 6.3250 1.0800 6.0050 1.0800 6.0050 0.6200 6.1250 0.6200
                 6.1250 0.9600 6.4450 0.9600 6.4450 1.0500 6.9850 1.0500 6.9850 0.6200 7.1050 0.6200
                 7.1050 1.3100 8.1450 1.3100 ;
        POLYGON  7.5250 0.8600 7.4050 0.8600 7.4050 0.6200 7.2250 0.6200 7.2250 0.5000 6.7450 0.5000
                 6.7450 0.8000 6.5050 0.8000 6.5050 0.6800 6.6250 0.6800 6.6250 0.3800 7.3450 0.3800
                 7.3450 0.5000 7.5250 0.5000 ;
        POLYGON  6.7650 2.1700 4.9100 2.1700 4.9100 2.0000 4.2350 2.0000 4.2350 2.2500 4.1150 2.2500
                 4.1150 2.0000 3.0150 2.0000 3.0150 2.0500 2.3850 2.0500 2.3850 2.0850 2.2650 2.0850
                 2.2650 1.8450 2.3700 1.8450 2.3700 1.1300 2.2650 1.1300 2.2650 0.6500 2.3850 0.6500
                 2.3850 1.0100 2.4900 1.0100 2.4900 1.9300 2.8950 1.9300 2.8950 1.8800 5.0300 1.8800
                 5.0300 2.0500 6.7650 2.0500 ;
        POLYGON  6.2050 1.3200 5.7650 1.3200 5.7650 0.4800 5.3250 0.4800 5.3250 0.3600 5.8850 0.3600
                 5.8850 1.2000 6.2050 1.2000 ;
        POLYGON  5.7250 1.6400 5.4850 1.6400 5.4850 1.5200 5.5250 1.5200 5.5250 1.2800 4.1150 1.2800
                 4.1150 1.1100 3.0950 1.1100 3.0950 1.1400 2.8550 1.1400 2.8550 1.0200 2.9750 1.0200
                 2.9750 0.9900 4.2350 0.9900 4.2350 1.1600 5.5250 1.1600 5.5250 0.6200 5.6450 0.6200
                 5.6450 1.5200 5.7250 1.5200 ;
        POLYGON  5.2250 0.8600 5.1350 0.8600 5.1350 1.0400 4.3550 1.0400 4.3550 0.8000 4.2350 0.8000
                 4.2350 0.6800 4.4750 0.6800 4.4750 0.9200 5.0150 0.9200 5.0150 0.7400 5.1050 0.7400
                 5.1050 0.6200 5.2250 0.6200 ;
        RECT  3.5550 1.6400 5.1250 1.7600 ;
        POLYGON  4.8950 0.8000 4.6550 0.8000 4.6550 0.5600 4.1150 0.5600 4.1150 0.7200 3.7950 0.7200
                 3.7950 0.8000 3.5550 0.8000 3.5550 0.6800 3.6750 0.6800 3.6750 0.6000 3.9950 0.6000
                 3.9950 0.4400 4.7750 0.4400 4.7750 0.6800 4.8950 0.6800 ;
        POLYGON  3.8750 0.4800 3.5550 0.4800 3.5550 0.5600 2.7750 0.5600 2.7750 0.8600 2.7350 0.8600
                 2.7350 1.5700 2.7750 1.5700 2.7750 1.8100 2.6550 1.8100 2.6550 1.6900 2.6150 1.6900
                 2.6150 0.7400 2.6550 0.7400 2.6550 0.5600 2.5550 0.5600 2.5550 0.5300 2.1450 0.5300
                 2.1450 1.1300 1.8050 1.1300 1.8050 1.2000 1.5650 1.2000 1.5650 1.0100 2.0250 1.0100
                 2.0250 0.4100 2.6750 0.4100 2.6750 0.4400 3.4350 0.4400 3.4350 0.3600 3.8750 0.3600 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END SDFFSRX1

MACRO SDFFSRHQX8
    CLASS CORE ;
    FOREIGN SDFFSRHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 16.2400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 1.3200 2.7750 2.1850 ;
        RECT  2.6550 0.6800 2.7750 0.9600 ;
        RECT  0.0700 1.2000 2.7550 1.3200 ;
        RECT  2.6350 0.8400 2.7550 1.4400 ;
        RECT  1.8150 0.6800 1.9350 2.1850 ;
        RECT  0.9750 0.6800 1.0950 2.1800 ;
        RECT  0.1350 0.6800 0.2550 2.1800 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 1.1700 5.2450 1.3900 ;
        RECT  4.9450 1.1700 5.2050 1.4100 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0950 2.1300 10.3150 2.2500 ;
        RECT  9.0950 1.7000 9.2150 2.2500 ;
        RECT  8.4950 1.7000 9.2150 1.8200 ;
        RECT  7.5350 2.1300 8.6150 2.2500 ;
        RECT  8.4950 1.7000 8.6150 2.2500 ;
        RECT  7.2950 2.0800 7.6550 2.2000 ;
        RECT  7.2950 1.4200 7.4150 2.2000 ;
        RECT  5.6100 1.4200 7.4150 1.5400 ;
        RECT  5.5800 1.2100 5.8050 1.4350 ;
        RECT  5.5800 1.1750 5.7300 1.4350 ;
        RECT  5.5650 1.2100 5.8050 1.3300 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.4150 0.9600 13.5350 1.2000 ;
        RECT  13.0650 0.9600 13.5350 1.0900 ;
        RECT  13.0650 0.9400 13.3250 1.0900 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.7550 0.7550 13.8750 1.1800 ;
        RECT  13.7000 1.0350 13.8500 1.4400 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  14.9350 1.2200 15.3550 1.4400 ;
        RECT  15.0950 1.2000 15.3550 1.4400 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  15.7300 1.1750 15.8800 1.4350 ;
        RECT  15.5550 0.9600 15.8500 1.2000 ;
        RECT  14.2350 0.9600 15.8500 1.0800 ;
        RECT  14.7350 0.9600 14.9750 1.1000 ;
        RECT  14.2350 0.9600 14.3550 1.4400 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 16.2400 0.1800 ;
        RECT  15.2950 -0.1800 15.4150 0.8400 ;
        RECT  13.7750 -0.1800 14.0150 0.3200 ;
        RECT  12.7250 -0.1800 12.9650 0.3200 ;
        RECT  10.6150 -0.1800 10.7350 0.6800 ;
        RECT  5.2650 0.6900 5.5050 0.8100 ;
        RECT  5.3850 -0.1800 5.5050 0.8100 ;
        RECT  3.9150 -0.1800 4.0350 0.6650 ;
        RECT  3.0750 -0.1800 3.1950 0.6650 ;
        RECT  2.2350 -0.1800 2.3550 0.6700 ;
        RECT  1.3950 -0.1800 1.5150 0.6700 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 16.2400 2.7900 ;
        RECT  15.0750 1.8000 15.1950 2.7900 ;
        RECT  13.7550 1.5600 13.8750 2.7900 ;
        RECT  12.8450 1.5600 12.9650 2.7900 ;
        RECT  10.4750 1.8800 10.7150 2.0000 ;
        RECT  10.4750 1.8800 10.5950 2.7900 ;
        RECT  8.8550 1.9400 8.9750 2.7900 ;
        RECT  8.7350 1.9400 8.9750 2.0600 ;
        RECT  6.6050 1.9000 6.8450 2.0200 ;
        RECT  6.6050 1.9000 6.7250 2.7900 ;
        RECT  5.2050 1.9000 5.4450 2.0200 ;
        RECT  5.2050 1.9000 5.3250 2.7900 ;
        RECT  3.9150 1.5350 4.0350 2.7900 ;
        RECT  3.0750 1.5350 3.1950 2.7900 ;
        RECT  2.2350 1.4400 2.3550 2.7900 ;
        RECT  1.3950 1.4400 1.5150 2.7900 ;
        RECT  0.5550 1.4400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  16.1200 1.9800 15.4350 1.9800 15.4350 1.8600 16.0000 1.8600 16.0000 1.6800
                 14.6350 1.6800 14.6350 1.4200 14.5150 1.4200 14.5150 1.3000 14.7550 1.3000
                 14.7550 1.5600 16.0000 1.5600 16.0000 0.8400 15.7150 0.8400 15.7150 0.6000
                 15.8350 0.6000 15.8350 0.7200 16.1200 0.7200 ;
        POLYGON  14.7150 0.6350 14.1150 0.6350 14.1150 1.5600 14.5150 1.5600 14.5150 2.2100
                 14.3950 2.2100 14.3950 1.6800 13.9950 1.6800 13.9950 0.6350 13.7300 0.6350
                 13.7300 0.5600 11.7950 0.5600 11.7950 1.0000 12.1350 1.0000 12.1350 1.5800
                 12.1550 1.5800 12.1550 1.7700 11.9150 1.7700 11.9150 1.5800 12.0150 1.5800
                 12.0150 1.1200 11.6750 1.1200 11.6750 0.4400 13.8500 0.4400 13.8500 0.5150
                 14.7150 0.5150 ;
        POLYGON  13.5150 1.7400 13.2750 1.7400 13.2750 1.4400 12.7250 1.4400 12.7250 2.2500
                 10.8350 2.2500 10.8350 1.7600 10.3550 1.7600 10.3550 2.0100 9.3350 2.0100
                 9.3350 1.5800 8.3750 1.5800 8.3750 2.0100 7.7750 2.0100 7.7750 0.9800 7.8750 0.9800
                 7.8750 0.4800 7.3950 0.4800 7.3950 1.0600 7.1550 1.0600 7.1550 0.9400 7.2750 0.9400
                 7.2750 0.3600 7.9950 0.3600 7.9950 1.1000 7.8950 1.1000 7.8950 1.8900 8.2550 1.8900
                 8.2550 1.4600 9.4550 1.4600 9.4550 1.8900 10.2350 1.8900 10.2350 1.6400 10.9550 1.6400
                 10.9550 2.1300 12.6050 2.1300 12.6050 0.7000 13.1950 0.7000 13.1950 0.6800
                 13.4350 0.6800 13.4350 0.8000 13.3150 0.8000 13.3150 0.8200 12.7250 0.8200
                 12.7250 1.3200 13.3950 1.3200 13.3950 1.6200 13.5150 1.6200 ;
        POLYGON  12.4850 2.0100 11.0750 2.0100 11.0750 1.2800 11.0550 1.2800 11.0550 1.1600
                 10.5750 1.1600 10.5750 1.2800 9.8150 1.2800 9.8150 1.1000 8.4750 1.1000 8.4750 1.0400
                 8.3550 1.0400 8.3550 0.9200 8.5950 0.9200 8.5950 0.9800 9.9350 0.9800 9.9350 1.1600
                 10.4550 1.1600 10.4550 1.0400 11.2950 1.0400 11.2950 1.1600 11.1950 1.1600
                 11.1950 1.8900 11.6750 1.8900 11.6750 1.3600 11.6550 1.3600 11.6550 1.2400
                 11.8950 1.2400 11.8950 1.3600 11.7950 1.3600 11.7950 1.8900 12.3650 1.8900
                 12.3650 0.8000 12.2450 0.8000 12.2450 0.6800 12.4850 0.6800 ;
        POLYGON  11.5550 1.7700 11.3150 1.7700 11.3150 1.6000 11.4150 1.6000 11.4150 0.7800
                 11.1100 0.7800 11.1100 0.9200 10.2950 0.9200 10.2950 1.0400 10.0550 1.0400
                 10.0550 0.9200 10.1750 0.9200 10.1750 0.8000 10.9900 0.8000 10.9900 0.6600
                 11.2550 0.6600 11.2550 0.5400 11.3750 0.5400 11.3750 0.6600 11.5350 0.6600
                 11.5350 1.6000 11.5550 1.6000 ;
        POLYGON  10.9350 1.4000 10.8150 1.4000 10.8150 1.5200 10.1150 1.5200 10.1150 1.7700
                 9.9950 1.7700 9.9950 1.5200 9.5750 1.5200 9.5750 1.3400 8.1350 1.3400 8.1350 1.7700
                 8.0150 1.7700 8.0150 1.2200 8.1150 1.2200 8.1150 0.5400 8.2350 0.5400 8.2350 0.6800
                 9.0400 0.6800 9.0400 0.7400 9.7150 0.7400 9.7150 0.6000 9.9550 0.6000 9.9550 0.7200
                 9.8350 0.7200 9.8350 0.8600 8.9200 0.8600 8.9200 0.8000 8.2350 0.8000 8.2350 1.2200
                 9.6950 1.2200 9.6950 1.4000 10.6950 1.4000 10.6950 1.2800 10.9350 1.2800 ;
        POLYGON  10.3150 0.6800 10.1950 0.6800 10.1950 0.4800 9.5350 0.4800 9.5350 0.6200 9.2950 0.6200
                 9.2950 0.5000 9.4150 0.5000 9.4150 0.3600 10.3150 0.3600 ;
        POLYGON  7.7550 0.7200 7.6550 0.7200 7.6550 1.9600 7.5350 1.9600 7.5350 1.3000 5.9250 1.3000
                 5.9250 1.0550 5.3650 1.0550 5.3650 1.0500 5.0250 1.0500 5.0250 0.4950 4.2750 0.4950
                 4.2750 1.1750 4.1550 1.1750 4.1550 0.3750 5.1450 0.3750 5.1450 0.9300 5.4850 0.9300
                 5.4850 0.9350 6.0450 0.9350 6.0450 1.1800 7.5350 1.1800 7.5350 0.7200 7.5150 0.7200
                 7.5150 0.6000 7.7550 0.6000 ;
        POLYGON  7.1750 1.9600 7.0550 1.9600 7.0550 1.7800 5.9250 1.7800 5.9250 1.9900 5.8050 1.9900
                 5.8050 1.6600 7.1750 1.6600 ;
        POLYGON  7.1550 0.7200 7.0350 0.7200 7.0350 1.0550 6.1650 1.0550 6.1650 0.6750 6.2850 0.6750
                 6.2850 0.9350 6.9150 0.9350 6.9150 0.6000 7.1550 0.6000 ;
        POLYGON  6.7050 0.8150 6.5850 0.8150 6.5850 0.5550 5.9100 0.5550 5.9100 0.5750 5.8650 0.5750
                 5.8650 0.8150 5.7450 0.8150 5.7450 0.4550 5.7900 0.4550 5.7900 0.4350 6.7050 0.4350 ;
        POLYGON  6.4850 2.2500 5.5650 2.2500 5.5650 1.7800 5.3000 1.7800 5.3000 1.7700 4.7850 1.7700
                 4.7850 1.6500 4.7050 1.6500 4.7050 0.9300 4.7850 0.9300 4.7850 0.6300 4.9050 0.6300
                 4.9050 1.0500 4.8250 1.0500 4.8250 1.5300 4.9050 1.5300 4.9050 1.6500 5.4200 1.6500
                 5.4200 1.6600 5.6850 1.6600 5.6850 2.1300 6.4850 2.1300 ;
        POLYGON  5.0850 2.2500 4.3350 2.2500 4.3350 1.5350 4.3950 1.5350 4.3950 1.4150 3.6150 1.4150
                 3.6150 2.1850 3.4950 2.1850 3.4950 1.2000 2.8750 1.2000 2.8750 1.0800 3.4950 1.0800
                 3.4950 0.6150 3.6150 0.6150 3.6150 1.2950 4.3950 1.2950 4.3950 0.6150 4.5150 0.6150
                 4.5150 1.6550 4.4550 1.6550 4.4550 2.1300 5.0850 2.1300 ;
    END
END SDFFSRHQX8

MACRO SDFFSRHQX4
    CLASS CORE ;
    FOREIGN SDFFSRHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.5000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.4450 1.5150 2.0950 ;
        RECT  1.3950 0.6300 1.5150 0.9700 ;
        RECT  1.3750 0.8500 1.4950 1.5650 ;
        RECT  0.5550 0.9700 1.4950 1.0900 ;
        RECT  0.5550 0.9400 0.8550 1.0900 ;
        RECT  0.5550 0.6300 0.6750 2.0950 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.0050 3.1200 1.4550 ;
        RECT  2.9700 0.9800 3.0900 1.4550 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.4300 1.2650 11.5500 1.5150 ;
        RECT  11.0350 1.2650 11.5500 1.3850 ;
        RECT  11.0350 1.2300 11.2950 1.3850 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6700 1.2800 12.0150 1.4850 ;
        RECT  11.6700 1.0900 11.8200 1.4850 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.3150 1.2350 13.6150 1.4650 ;
        RECT  13.3550 1.2100 13.6150 1.4650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.9850 0.9700 14.1050 1.2200 ;
        RECT  12.7350 0.9700 14.1050 1.0900 ;
        RECT  13.6450 0.9400 13.9050 1.0900 ;
        RECT  12.7350 0.9700 12.9750 1.1000 ;
        END
    END SE
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.3150 2.1300 8.5550 2.2500 ;
        RECT  7.6750 2.0100 8.4350 2.1300 ;
        RECT  7.6750 1.7000 7.7950 2.1300 ;
        RECT  7.0750 1.7000 7.7950 1.8200 ;
        RECT  5.7550 2.1300 7.1950 2.2500 ;
        RECT  7.0750 1.7000 7.1950 2.2500 ;
        RECT  5.7550 1.5200 5.8750 2.2500 ;
        RECT  5.2350 1.5200 5.8750 1.6400 ;
        RECT  5.2350 1.5200 5.4950 1.6700 ;
        RECT  5.0550 1.4700 5.3550 1.5900 ;
        END
    END SN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.5000 0.1800 ;
        RECT  14.2450 -0.1800 14.3650 0.8800 ;
        RECT  13.2350 0.4600 13.4750 0.5800 ;
        RECT  13.2350 -0.1800 13.3550 0.5800 ;
        RECT  11.8150 -0.1800 12.0550 0.3400 ;
        RECT  11.1850 -0.1800 11.4250 0.3800 ;
        RECT  9.1350 0.4600 9.3750 0.5800 ;
        RECT  9.1350 -0.1800 9.2550 0.5800 ;
        RECT  5.2050 -0.1800 5.3250 0.4600 ;
        RECT  2.5950 0.5000 2.8350 0.6200 ;
        RECT  2.7150 -0.1800 2.8350 0.6200 ;
        RECT  1.8150 -0.1800 1.9350 0.6800 ;
        RECT  0.9750 -0.1800 1.0950 0.6800 ;
        RECT  0.1350 -0.1800 0.2550 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.5000 2.7900 ;
        RECT  14.2450 1.4600 14.3650 2.7900 ;
        RECT  13.5150 1.8250 13.6350 2.7900 ;
        RECT  12.2350 1.7600 12.3550 2.7900 ;
        RECT  10.9750 1.9400 11.0950 2.7900 ;
        RECT  8.6750 2.0100 8.9150 2.1300 ;
        RECT  8.6750 2.0100 8.7950 2.7900 ;
        RECT  7.3150 1.9400 7.5550 2.0600 ;
        RECT  7.3150 1.9400 7.4350 2.7900 ;
        RECT  4.8550 2.2900 5.0950 2.7900 ;
        RECT  3.5950 2.1750 3.7150 2.7900 ;
        RECT  2.7150 2.1750 2.8350 2.7900 ;
        RECT  1.8150 1.5750 1.9350 2.7900 ;
        RECT  0.9750 1.4450 1.0950 2.7900 ;
        RECT  0.1350 1.4450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.0050 0.8200 13.3550 0.8200 13.3550 0.8500 12.6150 0.8500 12.6150 1.2200
                 13.1350 1.2200 13.1350 1.5850 13.7650 1.5850 13.7650 1.4950 14.0050 1.4950
                 14.0050 1.6150 13.8850 1.6150 13.8850 1.7050 13.0150 1.7050 13.0150 1.3400
                 12.4950 1.3400 12.4950 1.1000 12.3750 1.1000 12.3750 0.9800 12.4950 0.9800
                 12.4950 0.7300 13.2350 0.7300 13.2350 0.7000 14.0050 0.7000 ;
        POLYGON  12.9950 2.2100 12.8750 2.2100 12.8750 1.9450 12.7750 1.9450 12.7750 1.5800
                 12.1350 1.5800 12.1350 0.6100 11.7250 0.6100 11.7250 0.6200 10.9450 0.6200
                 10.9450 0.4800 10.3750 0.4800 10.3750 0.7200 10.1950 0.7200 10.1950 1.8000
                 10.1750 1.8000 10.1750 2.0100 10.0550 2.0100 10.0550 1.6800 10.0750 1.6800
                 10.0750 0.3600 11.0650 0.3600 11.0650 0.5000 11.6050 0.5000 11.6050 0.4900
                 12.7550 0.4900 12.7550 0.6100 12.2550 0.6100 12.2550 1.4600 12.8950 1.4600
                 12.8950 1.8250 12.9950 1.8250 ;
        POLYGON  11.9950 1.9400 11.4900 1.9400 11.4900 1.8200 10.6500 1.8200 10.6500 2.2500
                 9.3950 2.2500 9.3950 1.8900 7.9150 1.8900 7.9150 1.5800 6.9550 1.5800 6.9550 2.0100
                 6.2350 2.0100 6.2350 1.2900 6.2750 1.2900 6.2750 0.9100 6.3550 0.9100 6.3550 0.5500
                 5.8750 0.5500 5.8750 1.1100 5.6350 1.1100 5.6350 0.9900 5.7550 0.9900 5.7550 0.4300
                 6.4750 0.4300 6.4750 1.0300 6.3950 1.0300 6.3950 1.4100 6.3550 1.4100 6.3550 1.8900
                 6.8350 1.8900 6.8350 1.4600 8.0350 1.4600 8.0350 1.7700 9.3950 1.7700 9.3950 1.4200
                 9.6750 1.4200 9.6750 1.5400 9.5150 1.5400 9.5150 2.1300 10.5300 2.1300 10.5300 1.7000
                 10.7950 1.7000 10.7950 1.1000 10.7750 1.1000 10.7750 0.8600 11.4300 0.8600
                 11.4300 0.7400 11.6950 0.7400 11.6950 0.8600 11.5500 0.8600 11.5500 0.9800
                 10.9150 0.9800 10.9150 1.7000 11.6100 1.7000 11.6100 1.8200 11.9950 1.8200 ;
        POLYGON  10.8250 0.7200 10.6150 0.7200 10.6150 1.4600 10.6750 1.4600 10.6750 1.5800
                 10.4350 1.5800 10.4350 1.4600 10.4950 1.4600 10.4950 1.3200 10.3150 1.3200
                 10.3150 1.0800 10.4950 1.0800 10.4950 0.6000 10.8250 0.6000 ;
        POLYGON  9.9550 0.7400 9.9350 0.7400 9.9350 1.7800 9.7550 1.7800 9.7550 2.0100 9.6350 2.0100
                 9.6350 1.6600 9.8150 1.6600 9.8150 0.7400 9.6900 0.7400 9.6900 0.8200 8.8750 0.8200
                 8.8750 1.0000 8.6350 1.0000 8.6350 0.8800 8.7550 0.8800 8.7550 0.7000 9.5700 0.7000
                 9.5700 0.6200 9.8350 0.6200 9.8350 0.5000 9.9550 0.5000 ;
        POLYGON  9.6950 1.2400 8.3950 1.2400 8.3950 1.1000 6.8350 1.1000 6.8350 0.9800 8.5150 0.9800
                 8.5150 1.1200 9.4550 1.1200 9.4550 1.1000 9.6950 1.1000 ;
        POLYGON  9.2750 1.5400 8.4150 1.5400 8.4150 1.6500 8.1550 1.6500 8.1550 1.3400 6.7150 1.3400
                 6.7150 1.7700 6.4750 1.7700 6.4750 1.5300 6.5950 1.5300 6.5950 0.6000 6.7150 0.6000
                 6.7150 0.7400 7.9550 0.7400 7.9550 0.6000 8.1950 0.6000 8.1950 0.7200 8.0750 0.7200
                 8.0750 0.8600 6.7150 0.8600 6.7150 1.2200 8.2750 1.2200 8.2750 1.4200 9.2750 1.4200 ;
        POLYGON  8.5550 0.6800 8.4350 0.6800 8.4350 0.4800 7.8350 0.4800 7.8350 0.6200 7.5350 0.6200
                 7.5350 0.5000 7.7150 0.5000 7.7150 0.3600 8.5550 0.3600 ;
        POLYGON  6.2350 0.7900 6.1150 0.7900 6.1150 1.9900 5.9950 1.9900 5.9950 1.3500 4.8150 1.3500
                 4.8150 1.5700 4.3150 1.5700 4.3150 2.0100 3.6950 2.0100 3.6950 2.0550 2.5150 2.0550
                 2.5150 1.2550 2.6350 1.2550 2.6350 1.9350 3.5750 1.9350 3.5750 1.8900 4.1950 1.8900
                 4.1950 1.4500 4.6950 1.4500 4.6950 1.2300 5.9950 1.2300 5.9950 0.6700 6.2350 0.6700 ;
        POLYGON  5.6350 0.7900 5.3950 0.7900 5.3950 0.7000 4.9650 0.7000 4.9650 0.4800 4.4850 0.4800
                 4.4850 0.5000 4.4250 0.5000 4.4250 0.6200 4.1850 0.6200 4.1850 0.5000 4.3050 0.5000
                 4.3050 0.3800 4.3650 0.3800 4.3650 0.3600 5.0850 0.3600 5.0850 0.5800 5.5150 0.5800
                 5.5150 0.6700 5.6350 0.6700 ;
        POLYGON  5.6350 1.9300 4.4350 1.9300 4.4350 1.6900 4.5550 1.6900 4.5550 1.8100 5.3950 1.8100
                 5.3950 1.7900 5.6350 1.7900 ;
        POLYGON  5.6350 2.2500 5.2150 2.2500 5.2150 2.1700 4.6450 2.1700 4.6450 2.2500 3.8750 2.2500
                 3.8750 2.1300 4.5250 2.1300 4.5250 2.0500 5.3350 2.0500 5.3350 2.1300 5.6350 2.1300 ;
        POLYGON  4.8450 0.8600 4.5750 0.8600 4.5750 1.2800 3.7050 1.2800 3.7050 0.7200 3.5850 0.7200
                 3.5850 0.6000 3.8250 0.6000 3.8250 1.1600 4.4550 1.1600 4.4550 0.7400 4.6050 0.7400
                 4.6050 0.6000 4.8450 0.6000 ;
        POLYGON  4.3350 1.0400 4.0950 1.0400 4.0950 0.8600 3.9450 0.8600 3.9450 0.4800 3.0750 0.4800
                 3.0750 0.8600 2.3550 0.8600 2.3550 2.0950 2.2350 2.0950 2.2350 1.2100 1.6150 1.2100
                 1.6150 1.0900 2.2350 1.0900 2.2350 0.5400 2.3550 0.5400 2.3550 0.7400 2.9550 0.7400
                 2.9550 0.3600 4.0650 0.3600 4.0650 0.7400 4.2150 0.7400 4.2150 0.9200 4.3350 0.9200 ;
        POLYGON  3.5850 1.3300 3.3600 1.3300 3.3600 1.6950 3.3150 1.6950 3.3150 1.8150 3.1950 1.8150
                 3.1950 1.5750 3.2400 1.5750 3.2400 0.7200 3.1950 0.7200 3.1950 0.6000 3.4350 0.6000
                 3.4350 0.7200 3.3600 0.7200 3.3600 1.2100 3.5850 1.2100 ;
    END
END SDFFSRHQX4

MACRO SDFFSRHQX2
    CLASS CORE ;
    FOREIGN SDFFSRHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.3400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0800 1.0450 2.3200 1.2500 ;
        RECT  2.1000 1.0450 2.2500 1.4350 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.2700 2.1300 7.4700 2.2500 ;
        RECT  6.2700 1.7000 6.3900 2.2500 ;
        RECT  5.6700 1.7000 6.3900 1.8200 ;
        RECT  4.5900 2.1300 5.7900 2.2500 ;
        RECT  5.6700 1.7000 5.7900 2.2500 ;
        RECT  4.3500 2.0800 4.7100 2.2000 ;
        RECT  4.3500 1.4000 4.4700 2.2000 ;
        RECT  2.8800 1.4000 4.4700 1.5200 ;
        RECT  2.8800 1.2300 3.0000 1.5200 ;
        RECT  2.6800 1.1950 2.9200 1.3800 ;
        RECT  2.6250 1.2300 3.0000 1.3800 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5350 1.1600 10.6550 1.4000 ;
        RECT  10.1650 1.2300 10.6550 1.3800 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.8950 0.9400 11.0150 1.3050 ;
        RECT  10.8000 0.7850 10.9500 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 1.2300 12.4550 1.4300 ;
        RECT  12.0750 1.2450 12.4550 1.4200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.8300 1.1750 12.9800 1.4350 ;
        RECT  12.6950 0.9900 12.9500 1.2300 ;
        RECT  11.3750 0.9900 12.9500 1.1100 ;
        RECT  11.8750 0.9800 12.1150 1.1100 ;
        RECT  11.3750 0.9900 11.4950 1.4400 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6300 1.7550 0.8000 2.0150 ;
        RECT  0.6300 1.5400 0.7700 2.0150 ;
        RECT  0.6300 1.5400 0.7500 2.1900 ;
        RECT  0.5900 0.8000 0.7100 1.6600 ;
        RECT  0.5700 0.6800 0.6900 0.9200 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.3400 0.1800 ;
        RECT  12.4350 -0.1800 12.5550 0.8400 ;
        RECT  10.9150 -0.1800 11.1550 0.3200 ;
        RECT  9.9400 -0.1800 10.1800 0.3200 ;
        RECT  7.7900 -0.1800 7.9100 0.6400 ;
        RECT  2.4000 -0.1800 2.5200 0.6850 ;
        RECT  0.9900 -0.1800 1.1100 0.7400 ;
        RECT  0.1500 -0.1800 0.2700 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.3400 2.7900 ;
        RECT  12.2150 1.7950 12.3350 2.7900 ;
        RECT  10.8950 1.5600 11.0150 2.7900 ;
        RECT  10.0000 1.7600 10.1200 2.7900 ;
        RECT  7.6300 1.8800 7.8700 2.0000 ;
        RECT  7.6300 1.8800 7.7500 2.7900 ;
        RECT  6.0300 1.9400 6.1500 2.7900 ;
        RECT  5.9100 1.9400 6.1500 2.0600 ;
        RECT  3.6600 1.8800 3.9000 2.0000 ;
        RECT  3.6800 1.8800 3.8000 2.7900 ;
        RECT  2.4000 1.7950 2.5200 2.7900 ;
        RECT  2.2800 1.7950 2.5200 1.9150 ;
        RECT  1.0500 1.5400 1.1700 2.7900 ;
        RECT  0.2100 1.5400 0.3300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.2200 1.9750 12.5750 1.9750 12.5750 1.8550 13.1000 1.8550 13.1000 1.6750
                 11.8350 1.6750 11.8350 1.4200 11.6550 1.4200 11.6550 1.3000 11.9550 1.3000
                 11.9550 1.5550 13.1000 1.5550 13.1000 0.8700 12.8550 0.8700 12.8550 0.6000
                 12.9750 0.6000 12.9750 0.7500 13.2200 0.7500 ;
        POLYGON  11.8550 0.6650 11.2550 0.6650 11.2550 1.5600 11.6550 1.5600 11.6550 2.2100
                 11.5350 2.2100 11.5350 1.6800 11.1350 1.6800 11.1350 0.6650 10.8700 0.6650
                 10.8700 0.5600 8.9700 0.5600 8.9700 0.9000 9.2100 0.9000 9.2100 1.5400 9.3100 1.5400
                 9.3100 1.7700 9.0700 1.7700 9.0700 1.5400 9.0900 1.5400 9.0900 1.0200 8.8500 1.0200
                 8.8500 0.4400 10.9900 0.4400 10.9900 0.5450 11.8550 0.5450 ;
        POLYGON  10.6550 1.7400 10.4150 1.7400 10.4150 1.6400 9.8800 1.6400 9.8800 2.2500 7.9900 2.2500
                 7.9900 1.7600 7.5100 1.7600 7.5100 2.0100 6.5100 2.0100 6.5100 1.5800 5.5500 1.5800
                 5.5500 2.0100 4.8300 2.0100 4.8300 1.2600 4.8500 1.2600 4.8500 0.8400 4.9500 0.8400
                 4.9500 0.4800 4.4700 0.4800 4.4700 1.0400 4.2300 1.0400 4.2300 0.9200 4.3500 0.9200
                 4.3500 0.3600 5.0700 0.3600 5.0700 0.9600 4.9700 0.9600 4.9700 1.3800 4.9500 1.3800
                 4.9500 1.8900 5.4300 1.8900 5.4300 1.4600 6.6300 1.4600 6.6300 1.8900 7.3900 1.8900
                 7.3900 1.6400 8.1100 1.6400 8.1100 2.1300 9.7600 2.1300 9.7600 1.5200 9.8000 1.5200
                 9.8000 0.9200 10.3350 0.9200 10.3350 0.6800 10.5750 0.6800 10.5750 0.8000
                 10.4550 0.8000 10.4550 1.0400 9.9200 1.0400 9.9200 1.5200 10.5350 1.5200
                 10.5350 1.6200 10.6550 1.6200 ;
        POLYGON  9.7000 0.8000 9.6400 0.8000 9.6400 2.0100 8.2300 2.0100 8.2300 1.1600 7.7500 1.1600
                 7.7500 1.2800 6.9900 1.2800 6.9900 1.1000 5.5500 1.1000 5.5500 1.0400 5.4300 1.0400
                 5.4300 0.9200 5.6700 0.9200 5.6700 0.9800 7.1100 0.9800 7.1100 1.1600 7.6300 1.1600
                 7.6300 1.0400 8.2300 1.0400 8.2300 1.0000 8.4700 1.0000 8.4700 1.1200 8.3500 1.1200
                 8.3500 1.8900 8.8300 1.8900 8.8300 1.1400 8.9700 1.1400 8.9700 1.3800 8.9500 1.3800
                 8.9500 1.8900 9.5200 1.8900 9.5200 0.8000 9.4600 0.8000 9.4600 0.6800 9.7000 0.6800 ;
        POLYGON  8.7100 1.7700 8.4700 1.7700 8.4700 1.6000 8.5900 1.6000 8.5900 0.7400 8.2850 0.7400
                 8.2850 0.8800 7.7550 0.8800 7.7550 0.9200 7.4700 0.9200 7.4700 1.0400 7.2300 1.0400
                 7.2300 0.9200 7.3500 0.9200 7.3500 0.8000 7.6350 0.8000 7.6350 0.7600 8.1650 0.7600
                 8.1650 0.6200 8.4300 0.6200 8.4300 0.5000 8.5500 0.5000 8.5500 0.6200 8.7100 0.6200 ;
        POLYGON  8.1100 1.4000 7.9900 1.4000 7.9900 1.5200 7.2700 1.5200 7.2700 1.7700 7.1500 1.7700
                 7.1500 1.5200 6.7500 1.5200 6.7500 1.3400 5.3100 1.3400 5.3100 1.7700 5.0700 1.7700
                 5.0700 1.5000 5.1900 1.5000 5.1900 0.5400 5.3100 0.5400 5.3100 0.6800 6.1550 0.6800
                 6.1550 0.7400 6.8300 0.7400 6.8300 0.6000 7.1300 0.6000 7.1300 0.7200 6.9500 0.7200
                 6.9500 0.8600 6.0350 0.8600 6.0350 0.8000 5.3100 0.8000 5.3100 1.2200 6.8700 1.2200
                 6.8700 1.4000 7.8700 1.4000 7.8700 1.2800 8.1100 1.2800 ;
        POLYGON  7.4900 0.6800 7.3700 0.6800 7.3700 0.4800 6.7100 0.4800 6.7100 0.6200 6.4700 0.6200
                 6.4700 0.5000 6.5900 0.5000 6.5900 0.3600 7.4900 0.3600 ;
        POLYGON  4.8300 0.7200 4.7100 0.7200 4.7100 1.9600 4.5900 1.9600 4.5900 1.2800 3.1200 1.2800
                 3.1200 1.0750 2.6900 1.0750 2.6900 0.9250 2.1600 0.9250 2.1600 0.4800 1.3500 0.4800
                 1.3500 1.1800 1.2300 1.1800 1.2300 0.3600 2.2800 0.3600 2.2800 0.8050 2.8100 0.8050
                 2.8100 0.9550 3.2400 0.9550 3.2400 1.1600 4.5900 1.1600 4.5900 0.6000 4.8300 0.6000 ;
        POLYGON  4.2300 0.7200 4.1100 0.7200 4.1100 0.9250 3.3600 0.9250 3.3600 0.7250 3.1800 0.7250
                 3.1800 0.6050 3.4800 0.6050 3.4800 0.8050 3.9900 0.8050 3.9900 0.6000 4.2300 0.6000 ;
        POLYGON  4.2300 1.9600 4.1100 1.9600 4.1100 1.7600 3.0000 1.7600 3.0000 1.9750 2.8800 1.9750
                 2.8800 1.6400 4.2300 1.6400 ;
        POLYGON  3.7800 0.6850 3.6600 0.6850 3.6600 0.4850 2.9400 0.4850 2.9400 0.6850 2.8200 0.6850
                 2.8200 0.3650 3.7800 0.3650 ;
        POLYGON  3.5600 2.2500 3.0550 2.2500 3.0550 2.2150 2.6400 2.2150 2.6400 1.6750 1.8600 1.6750
                 1.8600 1.5500 1.8400 1.5500 1.8400 0.7200 1.8000 0.7200 1.8000 0.6000 2.0400 0.6000
                 2.0400 0.7200 1.9600 0.7200 1.9600 1.4300 1.9800 1.4300 1.9800 1.5550 2.7600 1.5550
                 2.7600 2.0950 3.1750 2.0950 3.1750 2.1300 3.5600 2.1300 ;
        POLYGON  2.2800 2.2500 2.0400 2.2500 2.0400 2.1800 1.4700 2.1800 1.4700 1.4200 0.8300 1.4200
                 0.8300 1.1800 0.9500 1.1800 0.9500 1.3000 1.4700 1.3000 1.4700 0.6000 1.5900 0.6000
                 1.5900 2.0600 2.1600 2.0600 2.1600 2.1300 2.2800 2.1300 ;
    END
END SDFFSRHQX2

MACRO SDFFSRHQX1
    CLASS CORE ;
    FOREIGN SDFFSRHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.4700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1400 1.9600 1.4350 ;
        RECT  1.7050 1.1100 1.8250 1.3950 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7300 2.1300 6.5900 2.2500 ;
        RECT  5.7300 1.9600 5.8500 2.2500 ;
        RECT  5.6300 1.7000 5.7500 2.0800 ;
        RECT  5.0300 1.7000 5.7500 1.8200 ;
        RECT  4.0700 2.1300 5.1500 2.2500 ;
        RECT  5.0300 1.7000 5.1500 2.2500 ;
        RECT  3.8300 2.0800 4.1900 2.2000 ;
        RECT  3.8300 1.4000 3.9500 2.2000 ;
        RECT  2.4200 1.4000 3.9500 1.5200 ;
        RECT  2.2200 1.1750 2.5400 1.4350 ;
        RECT  2.2200 1.1400 2.3400 1.4350 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 0.9550 9.7000 1.1200 ;
        RECT  9.2950 0.9400 9.5550 1.1450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.8200 0.8300 10.1700 1.1200 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.2600 1.2300 11.5850 1.3800 ;
        RECT  11.2600 1.2150 11.5300 1.5350 ;
        RECT  11.3200 1.2100 11.5300 1.5350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6500 0.9900 11.8900 1.1100 ;
        RECT  10.5300 0.9700 11.8750 1.0900 ;
        RECT  11.6150 0.9400 11.8750 1.0900 ;
        RECT  10.5300 0.9700 10.6500 1.4400 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1900 1.2950 0.3100 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.4700 0.1800 ;
        RECT  11.5900 -0.1800 11.7100 0.8200 ;
        RECT  10.0700 -0.1800 10.3100 0.3200 ;
        RECT  8.8350 -0.1800 9.0750 0.3200 ;
        RECT  7.0100 0.4900 7.2500 0.6100 ;
        RECT  7.0100 -0.1800 7.1300 0.6100 ;
        RECT  1.7600 -0.1800 2.0000 0.3200 ;
        RECT  0.5550 -0.1800 0.6750 0.8200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.4700 2.7900 ;
        RECT  11.3700 1.8950 11.4900 2.7900 ;
        RECT  10.0500 1.8500 10.1700 2.7900 ;
        RECT  9.3200 1.5050 9.4400 2.7900 ;
        RECT  6.7100 2.0100 6.9500 2.1300 ;
        RECT  6.7100 2.0100 6.8300 2.7900 ;
        RECT  5.3900 1.9400 5.5100 2.7900 ;
        RECT  5.2700 1.9400 5.5100 2.0600 ;
        RECT  3.1400 1.8800 3.3800 2.0000 ;
        RECT  3.1600 1.8800 3.2800 2.7900 ;
        RECT  1.8800 1.7950 2.0000 2.7900 ;
        RECT  1.7600 1.7950 2.0000 1.9150 ;
        RECT  0.6100 1.6900 0.7300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.1900 0.7600 12.1300 0.7600 12.1300 1.8950 11.9100 1.8950 11.9100 2.0900
                 11.7900 2.0900 11.7900 1.7750 10.9300 1.7750 10.9300 1.4200 10.8100 1.4200
                 10.8100 1.3000 11.0500 1.3000 11.0500 1.6550 12.0100 1.6550 12.0100 0.7600
                 11.9500 0.7600 11.9500 0.6400 12.1900 0.6400 ;
        POLYGON  11.0100 0.6100 10.7700 0.6100 10.7700 0.5600 10.4100 0.5600 10.4100 1.5600
                 10.8100 1.5600 10.8100 2.2100 10.6900 2.2100 10.6900 1.6800 10.2900 1.6800
                 10.2900 0.5600 8.2500 0.5600 8.2500 1.0400 8.6100 1.0400 8.6100 1.6200 8.6300 1.6200
                 8.6300 1.7700 8.3900 1.7700 8.3900 1.6200 8.4900 1.6200 8.4900 1.1600 8.1300 1.1600
                 8.1300 0.4400 10.8900 0.4400 10.8900 0.4900 11.0100 0.4900 ;
        POLYGON  9.8100 2.0750 9.5700 2.0750 9.5700 1.3850 9.2000 1.3850 9.2000 2.2500 7.2950 2.2500
                 7.2950 1.8900 5.9700 1.8900 5.9700 1.8400 5.8700 1.8400 5.8700 1.5800 4.9100 1.5800
                 4.9100 2.0100 4.3100 2.0100 4.3100 0.9800 4.4300 0.9800 4.4300 0.4800 3.9500 0.4800
                 3.9500 1.0400 3.6900 1.0400 3.6900 0.9200 3.8300 0.9200 3.8300 0.3600 4.5500 0.3600
                 4.5500 1.1000 4.4300 1.1000 4.4300 1.8900 4.7900 1.8900 4.7900 1.4600 5.9900 1.4600
                 5.9900 1.7200 6.0900 1.7200 6.0900 1.7700 7.4150 1.7700 7.4150 2.1300 9.0800 2.1300
                 9.0800 1.3850 9.0550 1.3850 9.0550 1.2200 8.9900 1.2200 8.9900 0.6800 9.4650 0.6800
                 9.4650 0.8000 9.1750 0.8000 9.1750 1.2650 9.6900 1.2650 9.6900 1.9550 9.8100 1.9550 ;
        POLYGON  8.9600 2.0100 7.5500 2.0100 7.5500 1.0900 7.0700 1.0900 7.0700 1.2100 7.0000 1.2100
                 7.0000 1.3600 6.3500 1.3600 6.3500 1.1000 4.9100 1.1000 4.9100 0.9800 6.4700 0.9800
                 6.4700 1.2400 6.8800 1.2400 6.8800 1.0900 6.9500 1.0900 6.9500 0.9700 7.7700 0.9700
                 7.7700 1.0900 7.6700 1.0900 7.6700 1.8900 8.1500 1.8900 8.1500 1.4000 8.1300 1.4000
                 8.1300 1.2800 8.3700 1.2800 8.3700 1.4000 8.2700 1.4000 8.2700 1.8900 8.8400 1.8900
                 8.8400 1.6250 8.7500 1.6250 8.7500 0.8400 8.4600 0.8400 8.4600 0.7200 8.8700 0.7200
                 8.8700 1.5050 8.9600 1.5050 ;
        POLYGON  8.0300 1.7700 7.7900 1.7700 7.7900 1.6200 7.8900 1.6200 7.8900 0.7700 7.5650 0.7700
                 7.5650 0.8500 6.8300 0.8500 6.8300 0.9700 6.7100 0.9700 6.7100 1.1200 6.5900 1.1200
                 6.5900 0.8500 6.7100 0.8500 6.7100 0.7300 7.4450 0.7300 7.4450 0.6500 7.7100 0.6500
                 7.7100 0.5300 7.8300 0.5300 7.8300 0.6500 8.0100 0.6500 8.0100 1.6200 8.0300 1.6200 ;
        POLYGON  7.4300 1.3300 7.3100 1.3300 7.3100 1.6000 6.4500 1.6000 6.4500 1.6500 6.2100 1.6500
                 6.2100 1.6000 6.1100 1.6000 6.1100 1.3400 4.6700 1.3400 4.6700 1.7700 4.5500 1.7700
                 4.5500 1.2200 4.6700 1.2200 4.6700 0.5400 4.7900 0.5400 4.7900 0.7400 5.9900 0.7400
                 5.9900 0.6000 6.2300 0.6000 6.2300 0.7200 6.1100 0.7200 6.1100 0.8600 4.7900 0.8600
                 4.7900 1.2200 6.2300 1.2200 6.2300 1.4800 7.1900 1.4800 7.1900 1.2100 7.4300 1.2100 ;
        POLYGON  6.5900 0.6800 6.4700 0.6800 6.4700 0.4800 5.8700 0.4800 5.8700 0.6200 5.5700 0.6200
                 5.5700 0.5000 5.7500 0.5000 5.7500 0.3600 6.5900 0.3600 ;
        POLYGON  4.3100 0.7200 4.1900 0.7200 4.1900 1.9600 4.0700 1.9600 4.0700 1.2800 2.6600 1.2800
                 2.6600 1.0200 2.0600 1.0200 2.0600 0.6000 1.3250 0.6000 1.3250 0.5600 0.9150 0.5600
                 0.9150 1.2600 0.7950 1.2600 0.7950 0.4400 1.4450 0.4400 1.4450 0.4800 2.1800 0.4800
                 2.1800 0.9000 2.7800 0.9000 2.7800 1.1600 4.0700 1.1600 4.0700 0.6000 4.3100 0.6000 ;
        POLYGON  3.7100 0.7200 3.5700 0.7200 3.5700 1.0200 2.9000 1.0200 2.9000 0.7800 2.6600 0.7800
                 2.6600 0.6600 3.0200 0.6600 3.0200 0.9000 3.4500 0.9000 3.4500 0.6000 3.7100 0.6000 ;
        POLYGON  3.7100 1.9600 3.5900 1.9600 3.5900 1.7600 2.4800 1.7600 2.4800 1.9800 2.3600 1.9800
                 2.3600 1.6400 3.7100 1.6400 ;
        POLYGON  3.2600 0.7800 3.1400 0.7800 3.1400 0.5400 2.4200 0.5400 2.4200 0.7800 2.3000 0.7800
                 2.3000 0.4200 3.2600 0.4200 ;
        POLYGON  3.0400 2.2500 2.8000 2.2500 2.8000 2.2200 2.1200 2.2200 2.1200 1.6750 1.3400 1.6750
                 1.3400 0.7200 1.6050 0.7200 1.6050 0.8400 1.4600 0.8400 1.4600 1.5550 2.2400 1.5550
                 2.2400 2.1000 2.9200 2.1000 2.9200 2.1300 3.0400 2.1300 ;
        POLYGON  1.7600 2.2500 1.0300 2.2500 1.0300 1.8200 1.0350 1.8200 1.0350 1.5000 0.4550 1.5000
                 0.4550 1.2400 0.5750 1.2400 0.5750 1.3800 1.0350 1.3800 1.0350 0.6800 1.1550 0.6800
                 1.1550 1.9400 1.1500 1.9400 1.1500 2.1300 1.7600 2.1300 ;
    END
END SDFFSRHQX1

MACRO SDFFSHQX8
    CLASS CORE ;
    FOREIGN SDFFSHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.9200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0350 1.4300 7.2750 1.5500 ;
        RECT  7.0350 1.4300 7.1550 1.8800 ;
        RECT  6.4650 1.7600 7.1550 1.8800 ;
        RECT  4.8850 1.8800 6.5850 2.0000 ;
        RECT  4.8850 1.2400 5.0250 1.4800 ;
        RECT  4.8850 1.2400 5.0050 2.0000 ;
        RECT  4.6550 1.5200 5.0050 1.6700 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7450 1.5200 11.0050 1.6950 ;
        RECT  10.6750 1.4350 10.9150 1.5850 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0350 1.2000 11.4050 1.3900 ;
        RECT  11.0350 1.1850 11.2950 1.4000 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.7750 1.2200 13.0350 1.4500 ;
        RECT  12.6850 1.2200 13.0350 1.4250 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.4100 1.1750 13.5600 1.4350 ;
        RECT  13.4100 0.9800 13.5300 1.4350 ;
        RECT  12.1850 0.9800 13.5300 1.1000 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5194  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1300 1.3500 3.2550 1.4700 ;
        RECT  3.1350 0.6500 3.2550 1.4700 ;
        RECT  3.0750 1.3500 3.1950 1.5900 ;
        RECT  2.2350 0.6500 2.3550 2.0900 ;
        RECT  2.1000 1.1050 2.3550 1.4350 ;
        RECT  0.5550 1.1050 2.3550 1.2250 ;
        RECT  1.3950 0.6500 1.5150 2.0900 ;
        RECT  0.5550 0.6550 0.6750 2.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.9200 0.1800 ;
        RECT  13.6650 -0.1800 13.7850 0.4000 ;
        RECT  12.8050 -0.1800 12.9250 0.6200 ;
        RECT  11.3450 0.4600 11.5850 0.5800 ;
        RECT  11.4650 -0.1800 11.5850 0.5800 ;
        RECT  10.1450 0.4650 10.3850 0.5850 ;
        RECT  10.2650 -0.1800 10.3850 0.5850 ;
        RECT  8.0350 -0.1800 8.1550 0.7300 ;
        RECT  6.8550 -0.1800 6.9750 0.6800 ;
        RECT  4.7650 0.5200 5.0050 0.6400 ;
        RECT  4.7650 -0.1800 4.8850 0.6400 ;
        RECT  3.9850 -0.1800 4.1050 0.7000 ;
        RECT  2.6550 -0.1800 2.7750 0.6400 ;
        RECT  1.8150 -0.1800 1.9350 0.6400 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.9200 2.7900 ;
        RECT  13.6650 2.0150 13.7850 2.7900 ;
        RECT  12.9050 1.8850 13.0250 2.7900 ;
        RECT  11.2650 1.5600 11.3850 2.7900 ;
        RECT  10.0350 1.4600 10.1550 2.7900 ;
        RECT  7.9050 2.2300 8.1450 2.7900 ;
        RECT  6.9450 2.2400 7.1850 2.7900 ;
        RECT  5.6050 2.1200 5.8450 2.2400 ;
        RECT  5.6050 2.1200 5.7250 2.7900 ;
        RECT  4.6450 2.1200 4.8850 2.2400 ;
        RECT  4.6450 2.1200 4.7650 2.7900 ;
        RECT  3.8050 1.5600 3.9250 2.7900 ;
        RECT  2.6550 1.5900 2.7750 2.7900 ;
        RECT  1.8150 1.3500 1.9350 2.7900 ;
        RECT  0.9750 1.3450 1.0950 2.7900 ;
        RECT  0.1350 1.3450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.3950 1.6750 13.2750 1.6750 13.2750 1.6900 12.4050 1.6900 12.4050 1.3400
                 11.8850 1.3400 11.8850 1.3700 11.7650 1.3700 11.7650 1.1300 11.9450 1.1300
                 11.9450 0.7400 13.3750 0.7400 13.3750 0.8600 12.0650 0.8600 12.0650 1.2200
                 12.5250 1.2200 12.5250 1.5700 13.1550 1.5700 13.1550 1.5550 13.3950 1.5550 ;
        POLYGON  12.3850 2.2100 12.2650 2.2100 12.2650 1.9300 12.1650 1.9300 12.1650 1.8100
                 11.5250 1.8100 11.5250 0.8200 11.1050 0.8200 11.1050 0.5300 10.6250 0.5300
                 10.6250 0.8250 9.9050 0.8250 9.9050 0.4800 9.3350 0.4800 9.3350 0.6100 9.4250 0.6100
                 9.4250 1.8100 9.3450 1.8100 9.3450 2.0100 9.2250 2.0100 9.2250 1.6900 9.3050 1.6900
                 9.3050 0.7300 9.2150 0.7300 9.2150 0.3600 10.0250 0.3600 10.0250 0.7050 10.5050 0.7050
                 10.5050 0.4100 11.2250 0.4100 11.2250 0.7000 11.7050 0.7000 11.7050 0.5000
                 12.2250 0.5000 12.2250 0.6200 11.8250 0.6200 11.8250 0.8200 11.6450 0.8200
                 11.6450 1.6900 12.2850 1.6900 12.2850 1.8100 12.3850 1.8100 ;
        POLYGON  10.9850 1.0650 10.5550 1.0650 10.5550 1.8150 10.8450 1.8150 10.8450 2.0550
                 10.7250 2.0550 10.7250 1.9350 10.4350 1.9350 10.4350 1.0650 9.8250 1.0650
                 9.8250 0.9450 10.7450 0.9450 10.7450 0.6500 10.9850 0.6500 ;
        POLYGON  9.7850 0.7200 9.7050 0.7200 9.7050 1.4600 9.7350 1.4600 9.7350 2.2500 8.2950 2.2500
                 8.2950 2.1100 7.6200 2.1100 7.6200 2.1200 6.8250 2.1200 6.8250 2.2400 6.1150 2.2400
                 6.1150 2.1200 6.7050 2.1200 6.7050 2.0000 7.5000 2.0000 7.5000 1.9900 8.4150 1.9900
                 8.4150 2.1300 8.9850 2.1300 8.9850 1.3700 9.1050 1.3700 9.1050 2.1300 9.6150 2.1300
                 9.6150 1.5800 9.5850 1.5800 9.5850 0.7200 9.5450 0.7200 9.5450 0.6000 9.7850 0.6000 ;
        POLYGON  9.1850 1.1500 9.0650 1.1500 9.0650 0.9700 8.9750 0.9700 8.9750 0.5300 8.4950 0.5300
                 8.4950 0.8900 8.6050 0.8900 8.6050 1.3300 8.6250 1.3300 8.6250 1.5700 8.5050 1.5700
                 8.5050 1.4500 8.4850 1.4500 8.4850 1.0100 8.3750 1.0100 8.3750 0.9700 7.7950 0.9700
                 7.7950 0.4800 7.3150 0.4800 7.3150 0.9200 6.8250 0.9200 6.8250 1.0400 6.5850 1.0400
                 6.5850 0.5000 5.7650 0.5000 5.7650 0.9800 5.8450 0.9800 5.8450 1.2200 5.6450 1.2200
                 5.6450 0.3800 6.7050 0.3800 6.7050 0.8000 7.1950 0.8000 7.1950 0.3600 7.9150 0.3600
                 7.9150 0.8500 8.3750 0.8500 8.3750 0.4100 9.0950 0.4100 9.0950 0.8500 9.1850 0.8500 ;
        POLYGON  8.8650 1.8100 8.8250 1.8100 8.8250 2.0100 8.7050 2.0100 8.7050 1.8100 8.2450 1.8100
                 8.2450 1.5300 7.6850 1.5300 7.6850 1.4100 8.3650 1.4100 8.3650 1.6900 8.7450 1.6900
                 8.7450 1.2100 8.7350 1.2100 8.7350 0.7700 8.6150 0.7700 8.6150 0.6500 8.8550 0.6500
                 8.8550 1.0900 8.8650 1.0900 ;
        POLYGON  8.3650 1.2800 7.5450 1.2800 7.5450 1.7500 7.6650 1.7500 7.6650 1.8700 7.4250 1.8700
                 7.4250 1.2800 6.8750 1.2800 6.8750 1.6400 6.7550 1.6400 6.7550 1.2800 6.3050 1.2800
                 6.3050 0.6400 6.4250 0.6400 6.4250 1.1600 7.4350 1.1600 7.4350 0.6000 7.6750 0.6000
                 7.6750 0.7200 7.5550 0.7200 7.5550 1.1600 8.3650 1.1600 ;
        POLYGON  6.4550 1.6400 6.3350 1.6400 6.3350 1.5200 6.0650 1.5200 6.0650 1.4600 5.1450 1.4600
                 5.1450 1.1200 4.7050 1.1200 4.7050 1.1500 4.4650 1.1500 4.4650 1.0000 5.2650 1.0000
                 5.2650 1.3400 5.9650 1.3400 5.9650 0.8600 5.8850 0.8600 5.8850 0.6200 6.0050 0.6200
                 6.0050 0.7400 6.0850 0.7400 6.0850 1.3400 6.1850 1.3400 6.1850 1.4000 6.4550 1.4000 ;
        RECT  5.1250 1.6400 6.0950 1.7600 ;
        POLYGON  5.5050 1.2000 5.3850 1.2000 5.3850 0.8800 4.3450 0.8800 4.3450 2.2100 4.2250 2.2100
                 4.2250 0.9400 3.6850 0.9400 3.6850 1.8600 3.5050 1.8600 3.5050 2.2100 3.3850 2.2100
                 3.3850 1.7400 3.5650 1.7400 3.5650 0.9400 3.3750 0.9400 3.3750 0.5300 3.0150 0.5300
                 3.0150 1.2300 2.8950 1.2300 2.8950 0.4100 3.4950 0.4100 3.4950 0.6500 3.6850 0.6500
                 3.6850 0.8200 4.2250 0.8200 4.2250 0.7600 4.4050 0.7600 4.4050 0.6400 4.5250 0.6400
                 4.5250 0.7600 5.5050 0.7600 ;
    END
END SDFFSHQX8

MACRO SDFFSHQX4
    CLASS CORE ;
    FOREIGN SDFFSHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.3300 1.5150 2.0800 ;
        RECT  1.3950 0.6300 1.5150 0.9700 ;
        RECT  1.3750 0.8500 1.4950 1.4500 ;
        RECT  0.5550 0.9700 1.4950 1.0900 ;
        RECT  0.5550 0.8850 0.8000 1.1450 ;
        RECT  0.5550 0.6300 0.6750 2.0800 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2050 1.4000 5.4450 1.5200 ;
        RECT  5.2050 1.4000 5.3250 1.7600 ;
        RECT  4.6150 1.7200 5.2650 1.8400 ;
        RECT  5.1450 1.6400 5.3250 1.7600 ;
        RECT  4.0850 1.8900 4.7350 2.0100 ;
        RECT  4.6150 1.7200 4.7350 2.0100 ;
        RECT  4.0850 1.7000 4.2050 2.0100 ;
        RECT  3.3750 1.7000 4.2050 1.8200 ;
        RECT  2.7100 1.9900 3.4950 2.1100 ;
        RECT  3.3750 1.7000 3.4950 2.1100 ;
        RECT  2.6750 1.1700 2.9150 1.2900 ;
        RECT  2.7100 1.1700 2.8300 2.1100 ;
        RECT  2.6800 1.4650 2.8300 1.7250 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7150 1.2100 8.9750 1.4500 ;
        RECT  8.6450 1.1150 8.8850 1.3300 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5150 0.9400 9.6350 1.1800 ;
        RECT  9.0050 0.9400 9.6350 1.0600 ;
        RECT  9.0050 0.9400 9.2650 1.0900 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0350 1.2200 11.3100 1.4150 ;
        RECT  11.0350 1.2200 11.1650 1.5550 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.3550 0.9800 11.9100 1.1000 ;
        RECT  11.6700 0.8850 11.8200 1.1450 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.9250 -0.1800 12.0450 0.7650 ;
        RECT  10.9750 -0.1800 11.0950 0.6200 ;
        RECT  9.4950 0.4600 9.7350 0.5800 ;
        RECT  9.6150 -0.1800 9.7350 0.5800 ;
        RECT  8.2950 -0.1800 8.5350 0.3200 ;
        RECT  6.3050 -0.1800 6.4250 0.6800 ;
        RECT  5.1250 -0.1800 5.2450 0.7200 ;
        RECT  2.6550 0.4500 2.8950 0.5700 ;
        RECT  2.6550 -0.1800 2.7750 0.5700 ;
        RECT  1.8150 -0.1800 1.9350 0.6800 ;
        RECT  0.9750 -0.1800 1.0950 0.6800 ;
        RECT  0.1350 -0.1800 0.2550 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.9250 1.4750 12.0450 2.7900 ;
        RECT  11.1950 1.9150 11.3150 2.7900 ;
        RECT  9.6350 1.5600 9.7550 2.7900 ;
        RECT  8.1650 1.4600 8.2850 2.7900 ;
        RECT  6.0550 2.2000 6.2950 2.7900 ;
        RECT  5.0950 2.2000 5.3350 2.7900 ;
        RECT  3.6150 1.9400 3.7350 2.7900 ;
        RECT  2.7150 2.2300 2.8350 2.7900 ;
        RECT  1.8750 2.2300 1.9950 2.7900 ;
        RECT  0.9750 1.4300 1.0950 2.7900 ;
        RECT  0.1350 1.4300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6850 0.7050 11.5500 0.7050 11.5500 0.8600 10.2350 0.8600 10.2350 1.3000
                 10.8750 1.3000 10.8750 1.4200 10.2350 1.4200 10.2350 1.6750 11.4450 1.6750
                 11.4450 1.5350 11.6850 1.5350 11.6850 1.6550 11.5650 1.6550 11.5650 1.7950
                 10.1150 1.7950 10.1150 1.0900 9.9950 1.0900 9.9950 0.9700 10.1150 0.9700
                 10.1150 0.7400 11.4300 0.7400 11.4300 0.5850 11.6850 0.5850 ;
        POLYGON  10.6750 2.2100 10.5550 2.2100 10.5550 2.0350 9.8750 2.0350 9.8750 1.4400 9.7550 1.4400
                 9.7550 0.8200 9.2550 0.8200 9.2550 0.5300 8.7750 0.5300 8.7750 0.5600 7.6050 0.5600
                 7.6050 1.8400 7.5350 1.8400 7.5350 2.0100 7.2950 2.0100 7.2950 1.7200 7.4850 1.7200
                 7.4850 0.4400 8.6550 0.4400 8.6550 0.4100 9.3750 0.4100 9.3750 0.7000 9.8700 0.7000
                 9.8700 0.5000 10.3750 0.5000 10.3750 0.6200 9.9900 0.6200 9.9900 0.8200 9.8750 0.8200
                 9.8750 1.3200 9.9950 1.3200 9.9950 1.9150 10.6750 1.9150 ;
        POLYGON  9.1350 0.8000 8.5250 0.8000 8.5250 1.5700 9.1350 1.5700 9.1350 1.8100 9.0150 1.8100
                 9.0150 1.6900 8.4050 1.6900 8.4050 1.1200 7.9650 1.1200 7.9650 1.0000 8.4050 1.0000
                 8.4050 0.6800 8.8950 0.6800 8.8950 0.6500 9.1350 0.6500 ;
        POLYGON  8.0550 0.8000 7.8450 0.8000 7.8450 1.3400 7.8650 1.3400 7.8650 2.2500 6.4450 2.2500
                 6.4450 2.0800 4.9750 2.0800 4.9750 2.2500 4.1250 2.2500 4.1250 2.1300 4.8550 2.1300
                 4.8550 1.9600 6.5650 1.9600 6.5650 2.1300 7.0550 2.1300 7.0550 1.3400 7.1750 1.3400
                 7.1750 2.1300 7.7450 2.1300 7.7450 1.4600 7.7250 1.4600 7.7250 0.6800 8.0550 0.6800 ;
        POLYGON  7.3650 1.1000 7.2450 1.1000 7.2450 0.4800 6.6950 0.4800 6.6950 1.2800 6.4550 1.2800
                 6.4550 1.1600 6.5750 1.1600 6.5750 0.9200 6.0650 0.9200 6.0650 0.5200 5.4850 0.5200
                 5.4850 0.9600 4.7050 0.9600 4.7050 0.4800 3.6350 0.4800 3.6350 0.9400 3.7950 0.9400
                 3.7950 1.0600 3.5150 1.0600 3.5150 0.3600 4.8250 0.3600 4.8250 0.8400 5.3650 0.8400
                 5.3650 0.4000 6.1850 0.4000 6.1850 0.8000 6.5750 0.8000 6.5750 0.3600 7.3650 0.3600 ;
        POLYGON  7.1250 0.7200 6.9350 0.7200 6.9350 2.0100 6.8150 2.0100 6.8150 1.5200 5.9550 1.5200
                 5.9550 1.5600 5.8350 1.5600 5.8350 1.3200 5.9550 1.3200 5.9550 1.4000 6.8150 1.4000
                 6.8150 0.6000 7.1250 0.6000 ;
        POLYGON  6.3350 1.2000 5.7150 1.2000 5.7150 1.7200 5.8150 1.7200 5.8150 1.8400 5.5750 1.8400
                 5.5750 1.7200 5.5950 1.7200 5.5950 1.2000 4.8850 1.2000 4.8850 1.6000 4.7650 1.6000
                 4.7650 1.2000 4.4650 1.2000 4.4650 0.7200 4.1750 0.7200 4.1750 0.6000 4.5850 0.6000
                 4.5850 1.0800 5.8250 1.0800 5.8250 0.7600 5.7050 0.7600 5.7050 0.6400 5.9450 0.6400
                 5.9450 1.0800 6.3350 1.0800 ;
        POLYGON  4.4650 1.7700 4.3450 1.7700 4.3450 1.4400 4.2250 1.4400 4.2250 1.3400 3.0350 1.3400
                 3.0350 1.0500 2.3150 1.0500 2.3150 0.9300 3.1550 0.9300 3.1550 1.2200 3.9150 1.2200
                 3.9150 0.7200 3.7550 0.7200 3.7550 0.6000 4.0350 0.6000 4.0350 1.2200 4.3450 1.2200
                 4.3450 1.3200 4.4650 1.3200 ;
        POLYGON  4.1050 1.5800 3.2550 1.5800 3.2550 1.8700 3.1350 1.8700 3.1350 1.4600 4.1050 1.4600 ;
        POLYGON  3.3950 1.1000 3.2750 1.1000 3.2750 0.8100 2.1950 0.8100 2.1950 1.4300 2.3550 1.4300
                 2.3550 1.9500 2.2350 1.9500 2.2350 1.5500 2.0750 1.5500 2.0750 1.2100 1.6150 1.2100
                 1.6150 1.0900 2.0750 1.0900 2.0750 0.6600 2.2350 0.6600 2.2350 0.5400 2.3550 0.5400
                 2.3550 0.6900 3.3950 0.6900 ;
    END
END SDFFSHQX4

MACRO SDFFSHQX2
    CLASS CORE ;
    FOREIGN SDFFSHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0850 1.4300 4.3250 1.5500 ;
        RECT  3.1750 1.7600 4.2050 1.8800 ;
        RECT  4.0850 1.4300 4.2050 1.8800 ;
        RECT  3.1750 1.7600 3.2950 2.0100 ;
        RECT  2.8350 1.8900 3.2950 2.0100 ;
        RECT  1.8250 1.9900 2.9550 2.1100 ;
        RECT  1.7750 1.2300 2.0150 1.4700 ;
        RECT  1.8250 1.2300 1.9450 2.1100 ;
        RECT  1.7550 1.2300 2.0150 1.3800 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8450 1.4050 8.1550 1.6500 ;
        RECT  7.8450 1.4050 8.1050 1.6700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2750 1.0550 8.5150 1.2650 ;
        RECT  8.1350 0.9400 8.3950 1.1750 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.8550 1.2200 10.1350 1.4150 ;
        RECT  9.8550 1.2200 9.9750 1.5550 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5100 0.8850 10.6600 1.1450 ;
        RECT  10.5100 0.8850 10.6300 1.1650 ;
        RECT  9.2350 0.9800 10.6600 1.1000 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6800 0.6750 1.9900 ;
        RECT  0.3050 0.9400 0.6750 1.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.7450 -0.1800 10.8650 0.7650 ;
        RECT  9.8550 -0.1800 9.9750 0.6200 ;
        RECT  8.3750 0.4600 8.6150 0.5800 ;
        RECT  8.4950 -0.1800 8.6150 0.5800 ;
        RECT  7.1750 -0.1800 7.4150 0.3800 ;
        RECT  5.1850 -0.1800 5.3050 0.7500 ;
        RECT  4.0050 -0.1800 4.1250 0.6800 ;
        RECT  1.7550 0.5100 1.9950 0.6300 ;
        RECT  1.7550 -0.1800 1.8750 0.6300 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.7450 1.4750 10.8650 2.7900 ;
        RECT  10.0150 1.9150 10.1350 2.7900 ;
        RECT  8.5150 1.5600 8.6350 2.7900 ;
        RECT  7.1750 1.4600 7.2950 2.7900 ;
        RECT  4.8650 2.2300 5.1050 2.7900 ;
        RECT  3.9050 2.2400 4.1450 2.7900 ;
        RECT  2.5450 2.2300 2.7850 2.7900 ;
        RECT  1.5850 2.2300 1.8250 2.7900 ;
        RECT  0.9750 1.3400 1.0950 2.7900 ;
        RECT  0.1350 1.3400 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.5050 0.7050 10.3850 0.7050 10.3850 0.8600 9.1150 0.8600 9.1150 1.3000 9.7350 1.3000
                 9.7350 1.6750 10.2650 1.6750 10.2650 1.5350 10.5050 1.5350 10.5050 1.6550
                 10.3850 1.6550 10.3850 1.7950 9.6150 1.7950 9.6150 1.4200 8.9950 1.4200 8.9950 1.0900
                 8.8750 1.0900 8.8750 0.9700 8.9950 0.9700 8.9950 0.7400 10.2650 0.7400 10.2650 0.5850
                 10.5050 0.5850 ;
        POLYGON  9.4950 2.2100 9.3750 2.2100 9.3750 1.6600 8.7550 1.6600 8.7550 1.4400 8.6350 1.4400
                 8.6350 0.8200 8.1350 0.8200 8.1350 0.5300 7.6550 0.5300 7.6550 0.6200 6.4850 0.6200
                 6.4850 1.7500 6.5050 1.7500 6.5050 2.0100 6.2650 2.0100 6.2650 1.7500 6.3650 1.7500
                 6.3650 0.5000 7.5350 0.5000 7.5350 0.4100 8.2550 0.4100 8.2550 0.7000 8.7500 0.7000
                 8.7500 0.5000 9.2550 0.5000 9.2550 0.6200 8.8700 0.6200 8.8700 0.8200 8.7550 0.8200
                 8.7550 1.3200 8.8750 1.3200 8.8750 1.5400 9.4950 1.5400 ;
        POLYGON  8.0150 0.8600 7.7250 0.8600 7.7250 1.7900 7.9550 1.7900 7.9550 2.0300 7.8350 2.0300
                 7.8350 1.9100 7.6050 1.9100 7.6050 1.1900 6.9750 1.1900 6.9750 1.0700 7.6050 1.0700
                 7.6050 0.7400 7.7750 0.7400 7.7750 0.6500 8.0150 0.6500 ;
        POLYGON  6.9350 0.8600 6.8550 0.8600 6.8550 1.4600 6.8750 1.4600 6.8750 2.2500 5.4950 2.2500
                 5.4950 2.1100 4.5950 2.1100 4.5950 2.1200 3.5350 2.1200 3.5350 2.2500 3.0750 2.2500
                 3.0750 2.1300 3.4150 2.1300 3.4150 2.0000 4.4750 2.0000 4.4750 1.9900 5.6150 1.9900
                 5.6150 2.1300 6.0250 2.1300 6.0250 1.3700 6.1450 1.3700 6.1450 2.1300 6.7550 2.1300
                 6.7550 1.5800 6.7350 1.5800 6.7350 0.8600 6.6950 0.8600 6.6950 0.7400 6.9350 0.7400 ;
        POLYGON  6.2450 1.1700 6.1250 1.1700 6.1250 0.5500 5.6450 0.5500 5.6450 1.2700 5.6650 1.2700
                 5.6650 1.3900 5.4250 1.3900 5.4250 1.2700 5.5250 1.2700 5.5250 0.9900 4.9450 0.9900
                 4.9450 0.4800 4.4650 0.4800 4.4650 0.9200 3.8950 0.9200 3.8950 1.0400 3.6550 1.0400
                 3.6550 0.9200 3.6950 0.9200 3.6950 0.4800 2.7550 0.4800 2.7550 0.9600 2.8350 0.9600
                 2.8350 1.2000 2.6350 1.2000 2.6350 0.3600 3.8150 0.3600 3.8150 0.8000 4.3450 0.8000
                 4.3450 0.3600 5.0650 0.3600 5.0650 0.8700 5.5250 0.8700 5.5250 0.4300 6.2450 0.4300 ;
        POLYGON  6.0050 0.7900 5.9050 0.7900 5.9050 1.6300 5.8550 1.6300 5.8550 2.0100 5.7350 2.0100
                 5.7350 1.6300 4.7050 1.6300 4.7050 1.3500 4.8250 1.3500 4.8250 1.5100 5.7850 1.5100
                 5.7850 0.7900 5.7650 0.7900 5.7650 0.6700 6.0050 0.6700 ;
        POLYGON  5.3050 1.2300 4.5650 1.2300 4.5650 1.7500 4.6250 1.7500 4.6250 1.8700 4.3850 1.8700
                 4.3850 1.7500 4.4450 1.7500 4.4450 1.2300 4.1350 1.2300 4.1350 1.3100 3.8350 1.3100
                 3.8350 1.6400 3.7150 1.6400 3.7150 1.2800 3.4150 1.2800 3.4150 0.8400 3.2950 0.8400
                 3.2950 0.6000 3.4150 0.6000 3.4150 0.7200 3.5350 0.7200 3.5350 1.1600 4.0150 1.1600
                 4.0150 1.1100 4.5850 1.1100 4.5850 0.6000 4.8250 0.6000 4.8250 0.7200 4.7050 0.7200
                 4.7050 1.1100 5.3050 1.1100 ;
        POLYGON  3.4150 1.6400 3.2950 1.6400 3.2950 1.5200 3.1750 1.5200 3.1750 1.4400 2.1350 1.4400
                 2.1350 1.1100 1.4550 1.1100 1.4550 0.9900 2.2550 0.9900 2.2550 1.3200 2.9550 1.3200
                 2.9550 0.8400 2.8750 0.8400 2.8750 0.6000 2.9950 0.6000 2.9950 0.7200 3.0750 0.7200
                 3.0750 1.3200 3.2950 1.3200 3.2950 1.4000 3.4150 1.4000 ;
        POLYGON  3.0550 1.7700 2.3050 1.7700 2.3050 1.8700 2.0650 1.8700 2.0650 1.7500 2.1850 1.7500
                 2.1850 1.6500 2.8150 1.6500 2.8150 1.5600 3.0550 1.5600 ;
        POLYGON  2.4950 1.1600 2.3750 1.1600 2.3750 0.8700 1.3350 0.8700 1.3350 1.3400 1.5150 1.3400
                 1.5150 1.8600 1.3950 1.8600 1.3950 1.4600 1.2150 1.4600 1.2150 1.2000 0.7950 1.2000
                 0.7950 1.0800 1.2150 1.0800 1.2150 0.7100 1.3950 0.7100 1.3950 0.5900 1.5150 0.5900
                 1.5150 0.7500 2.4950 0.7500 ;
    END
END SDFFSHQX2

MACRO SDFFSHQX1
    CLASS CORE ;
    FOREIGN SDFFSHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.4300 4.0250 1.5500 ;
        RECT  2.8450 1.7500 3.9050 1.8700 ;
        RECT  3.7850 1.4300 3.9050 1.8700 ;
        RECT  2.8450 1.7500 2.9650 2.0100 ;
        RECT  2.3150 1.8900 2.9650 2.0100 ;
        RECT  1.5750 1.9900 2.4350 2.1100 ;
        RECT  1.5750 1.3500 1.7300 1.5900 ;
        RECT  1.5750 1.3500 1.6950 2.1100 ;
        RECT  1.5200 1.4650 1.6950 1.7250 ;
        END
    END SN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2450 1.2300 7.6100 1.3900 ;
        RECT  7.2450 1.2300 7.6050 1.4250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.4100 0.9400 7.8250 1.1100 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0050 1.2000 9.2650 1.4300 ;
        RECT  9.1050 1.2000 9.2250 1.6100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.7150 0.9600 9.8350 1.2000 ;
        RECT  9.6400 0.8850 9.7900 1.1450 ;
        RECT  8.4850 0.9600 9.8350 1.0800 ;
        RECT  8.4850 0.9600 8.7250 1.0900 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2696  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.6750 1.2200 1.0900 1.3400 ;
        RECT  0.6750 0.7200 0.9150 0.8400 ;
        RECT  0.6750 0.7200 0.7950 1.4600 ;
        RECT  0.6050 1.3400 0.7250 1.5800 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  9.9950 -0.1800 10.1150 0.7650 ;
        RECT  9.1050 -0.1800 9.2250 0.6000 ;
        RECT  7.6250 0.4600 7.8650 0.5800 ;
        RECT  7.7450 -0.1800 7.8650 0.5800 ;
        RECT  6.4250 -0.1800 6.6650 0.3400 ;
        RECT  4.8250 -0.1800 4.9450 0.7500 ;
        RECT  3.6450 -0.1800 3.7650 0.6500 ;
        RECT  1.5300 0.5000 1.7700 0.6200 ;
        RECT  1.5300 -0.1800 1.6500 0.6200 ;
        RECT  0.0750 0.5300 0.3150 0.6500 ;
        RECT  0.0750 -0.1800 0.1950 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  10.0550 1.9800 10.1750 2.7900 ;
        RECT  9.2650 1.9700 9.3850 2.7900 ;
        RECT  7.6850 1.5600 7.8050 2.7900 ;
        RECT  6.7550 1.4600 6.8750 2.7900 ;
        RECT  4.5950 2.2300 4.8350 2.7900 ;
        RECT  3.6350 2.2300 3.8750 2.7900 ;
        RECT  2.2950 2.2300 2.5350 2.7900 ;
        RECT  1.3350 2.2300 1.5750 2.7900 ;
        RECT  0.1850 1.3400 0.3050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.7550 0.7050 9.5200 0.7050 9.5200 0.8400 8.3650 0.8400 8.3650 1.2100 8.8850 1.2100
                 8.8850 1.7300 9.3450 1.7300 9.3450 1.5500 9.5150 1.5500 9.5150 1.5200 9.7550 1.5200
                 9.7550 1.6700 9.4650 1.6700 9.4650 1.8500 8.7650 1.8500 8.7650 1.3300 8.1850 1.3300
                 8.1850 0.9400 8.2450 0.9400 8.2450 0.7200 9.4000 0.7200 9.4000 0.5850 9.7550 0.5850 ;
        POLYGON  8.7450 2.2100 8.6250 2.2100 8.6250 2.0900 8.5250 2.0900 8.5250 1.5700 7.9450 1.5700
                 7.9450 0.8200 7.3850 0.8200 7.3850 0.5300 6.9050 0.5300 6.9050 0.5800 6.1550 0.5800
                 6.1550 1.7900 6.1750 1.7900 6.1750 2.0100 5.9350 2.0100 5.9350 1.7900 6.0350 1.7900
                 6.0350 0.8100 5.9450 0.8100 5.9450 0.4600 6.7850 0.4600 6.7850 0.4100 7.5050 0.4100
                 7.5050 0.7000 8.0000 0.7000 8.0000 0.4800 8.5050 0.4800 8.5050 0.6000 8.1200 0.6000
                 8.1200 0.8200 8.0650 0.8200 8.0650 1.4500 8.6450 1.4500 8.6450 1.9700 8.7450 1.9700 ;
        POLYGON  7.3250 1.8000 7.2050 1.8000 7.2050 1.6650 7.0050 1.6650 7.0050 1.1900 6.5550 1.1900
                 6.5550 1.0700 7.0050 1.0700 7.0050 0.7000 7.0250 0.7000 7.0250 0.6500 7.2650 0.6500
                 7.2650 0.8200 7.1250 0.8200 7.1250 1.5450 7.3250 1.5450 ;
        POLYGON  6.5150 0.8600 6.4350 0.8600 6.4350 1.3400 6.4550 1.3400 6.4550 2.2500 5.1650 2.2500
                 5.1650 2.1100 3.2050 2.1100 3.2050 2.2500 2.8050 2.2500 2.8050 2.1300 3.0850 2.1300
                 3.0850 1.9900 5.2850 1.9900 5.2850 2.1300 5.6950 2.1300 5.6950 1.3700 5.8150 1.3700
                 5.8150 2.1300 6.3350 2.1300 6.3350 1.4600 6.3150 1.4600 6.3150 0.8600 6.2750 0.8600
                 6.2750 0.7400 6.5150 0.7400 ;
        POLYGON  5.9150 1.1700 5.7950 1.1700 5.7950 1.0500 5.7050 1.0500 5.7050 0.4900 5.3350 0.4900
                 5.3350 1.5700 5.2150 1.5700 5.2150 0.9900 4.5850 0.9900 4.5850 0.4800 4.1750 0.4800
                 4.1750 0.8900 3.4900 0.8900 3.4900 0.9900 3.3700 0.9900 3.3700 0.4800 2.4500 0.4800
                 2.4500 0.8800 2.5500 0.8800 2.5500 1.1200 2.3300 1.1200 2.3300 0.3600 3.4900 0.3600
                 3.4900 0.7700 4.0550 0.7700 4.0550 0.3600 4.7050 0.3600 4.7050 0.8700 5.2150 0.8700
                 5.2150 0.3700 5.8250 0.3700 5.8250 0.9300 5.9150 0.9300 ;
        POLYGON  5.5850 0.8500 5.5750 0.8500 5.5750 1.8100 5.5350 1.8100 5.5350 2.0100 5.4150 2.0100
                 5.4150 1.8100 4.4750 1.8100 4.4750 1.5900 4.4350 1.5900 4.4350 1.3500 4.5550 1.3500
                 4.5550 1.4700 4.5950 1.4700 4.5950 1.6900 5.4550 1.6900 5.4550 0.7300 5.4650 0.7300
                 5.4650 0.6100 5.5850 0.6100 ;
        POLYGON  5.0550 1.2300 4.3150 1.2300 4.3150 1.7500 4.3550 1.7500 4.3550 1.8700 4.1150 1.8700
                 4.1150 1.7500 4.1950 1.7500 4.1950 1.2300 3.5650 1.2300 3.5650 1.6300 3.4450 1.6300
                 3.4450 1.2300 3.1300 1.2300 3.1300 0.7200 2.9900 0.7200 2.9900 0.6000 3.2500 0.6000
                 3.2500 1.1100 4.3450 1.1100 4.3450 0.6000 4.4650 0.6000 4.4650 1.1100 5.0550 1.1100 ;
        POLYGON  3.1450 1.6300 3.0250 1.6300 3.0250 1.4700 2.8900 1.4700 2.8900 1.3600 1.8500 1.3600
                 1.8500 1.1900 1.4500 1.1900 1.4500 1.0700 1.9700 1.0700 1.9700 1.2400 2.6700 1.2400
                 2.6700 0.7200 2.5700 0.7200 2.5700 0.6000 2.8100 0.6000 2.8100 0.7200 2.7900 0.7200
                 2.7900 1.2400 3.0100 1.2400 3.0100 1.3500 3.1450 1.3500 ;
        POLYGON  2.7250 1.7700 2.0550 1.7700 2.0550 1.8700 1.8150 1.8700 1.8150 1.7500 1.9350 1.7500
                 1.9350 1.6500 2.6050 1.6500 2.6050 1.4800 2.7250 1.4800 ;
        POLYGON  2.2100 1.1000 2.0900 1.1000 2.0900 0.8600 1.3300 0.8600 1.3300 1.6750 1.0350 1.6750
                 1.0350 2.2100 0.9150 2.2100 0.9150 1.5550 1.2100 1.5550 1.2100 0.8600 1.0350 0.8600
                 1.0350 0.6000 0.5550 0.6000 0.5550 1.2200 0.4350 1.2200 0.4350 0.4800 1.1550 0.4800
                 1.1550 0.5400 1.2900 0.5400 1.2900 0.6600 1.3300 0.6600 1.3300 0.7400 2.2100 0.7400 ;
    END
END SDFFSHQX1

MACRO SDFFRXL
    CLASS CORE ;
    FOREIGN SDFFRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4650 2.0950 1.6750 ;
        RECT  1.9750 1.3200 2.0950 1.6750 ;
        RECT  1.8100 1.4650 1.9600 1.8150 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3012  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 2.5100  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 1.2500 3.3350 1.4150 ;
        RECT  2.9150 1.2300 3.1750 1.4300 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0350 0.7600 8.1550 1.0300 ;
        RECT  7.9000 0.8600 8.0500 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 0.9600 9.5750 1.2000 ;
        RECT  9.2950 0.9400 9.5550 1.2000 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.8750 0.9400 10.1350 1.0900 ;
        RECT  9.7950 0.7000 9.9300 1.0600 ;
        RECT  8.6550 0.7000 9.9300 0.8200 ;
        RECT  9.0550 0.7000 9.1750 0.9800 ;
        RECT  8.5150 1.1000 8.7750 1.2200 ;
        RECT  8.6550 0.7000 8.7750 1.2200 ;
        RECT  8.5150 1.1000 8.6350 1.3400 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3350 1.4650 1.6700 1.7250 ;
        RECT  1.3750 0.6800 1.4950 0.9600 ;
        RECT  1.3350 0.8400 1.4550 2.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  9.4750 0.4600 9.7150 0.5800 ;
        RECT  9.4750 -0.1800 9.5950 0.5800 ;
        RECT  8.0350 -0.1800 8.1550 0.6400 ;
        RECT  5.3550 -0.1800 5.5950 0.3700 ;
        RECT  3.2950 0.4900 3.5350 0.6100 ;
        RECT  3.2950 -0.1800 3.4150 0.6100 ;
        RECT  1.7750 -0.1800 1.8950 0.4000 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  9.5350 1.5600 9.6550 2.7900 ;
        RECT  8.0950 2.0800 8.2150 2.7900 ;
        RECT  5.9950 2.1500 6.1150 2.7900 ;
        RECT  5.0950 2.2900 5.3350 2.7900 ;
        RECT  3.4650 2.2900 3.7050 2.7900 ;
        RECT  2.5650 2.0500 2.6850 2.7900 ;
        RECT  1.7550 1.9700 1.8750 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.3750 1.5600 10.0750 1.5600 10.0750 1.6800 9.9550 1.6800 9.9550 1.4400 9.0150 1.4400
                 9.0150 1.3000 8.8950 1.3000 8.8950 1.1800 9.1350 1.1800 9.1350 1.3200 10.2550 1.3200
                 10.2550 0.5800 9.8950 0.5800 9.8950 0.4600 10.3750 0.4600 ;
        POLYGON  9.0750 0.5800 8.5350 0.5800 8.5350 0.9800 8.3950 0.9800 8.3950 1.5000 8.8550 1.5000
                 8.8550 1.6200 8.3950 1.6200 8.3950 1.8600 7.2250 1.8600 7.2250 1.3600 6.8950 1.3600
                 6.8950 0.6200 7.0150 0.6200 7.0150 1.2400 7.3450 1.2400 7.3450 1.7400 8.2750 1.7400
                 8.2750 0.8600 8.4150 0.8600 8.4150 0.4600 9.0750 0.4600 ;
        POLYGON  7.9550 2.1000 6.6450 2.1000 6.6450 2.0800 6.3800 2.0800 6.3800 2.0300 5.8500 2.0300
                 5.8500 1.9300 2.3750 1.9300 2.3750 1.9700 2.2950 1.9700 2.2950 2.0900 2.1750 2.0900
                 2.1750 1.8100 2.2550 1.8100 2.2550 0.6800 2.3750 0.6800 2.3750 1.8100 3.8950 1.8100
                 3.8950 0.9700 4.0350 0.9700 4.0350 1.2100 4.0150 1.2100 4.0150 1.8100 4.4950 1.8100
                 4.4950 1.3700 4.4350 1.3700 4.4350 1.2500 4.6750 1.2500 4.6750 1.3700 4.6150 1.3700
                 4.6150 1.8100 5.9700 1.8100 5.9700 1.9100 6.5000 1.9100 6.5000 1.9600 6.6450 1.9600
                 6.6450 1.8400 6.7650 1.8400 6.7650 1.9800 7.9550 1.9800 ;
        POLYGON  7.7950 1.6200 7.5550 1.6200 7.5550 1.0000 7.3550 1.0000 7.3550 1.1200 7.2350 1.1200
                 7.2350 0.5000 6.2950 0.5000 6.2950 0.6100 5.1150 0.6100 5.1150 0.5600 4.6350 0.5600
                 4.6350 0.9700 4.9750 0.9700 4.9750 1.2100 4.8550 1.2100 4.8550 1.0900 4.5150 1.0900
                 4.5150 0.4400 5.2350 0.4400 5.2350 0.4900 6.1750 0.4900 6.1750 0.3600 6.4150 0.3600
                 6.4150 0.3800 7.3550 0.3800 7.3550 0.8800 7.5550 0.8800 7.5550 0.4000 7.6750 0.4000
                 7.6750 1.5000 7.7950 1.5000 ;
        POLYGON  6.9250 1.7200 6.8050 1.7200 6.8050 1.6000 6.6250 1.6000 6.6250 1.3600 5.3350 1.3600
                 5.3350 0.9700 5.4550 0.9700 5.4550 1.2400 6.4750 1.2400 6.4750 0.6200 6.5950 0.6200
                 6.5950 1.2400 6.7450 1.2400 6.7450 1.4800 6.9250 1.4800 ;
        POLYGON  6.5050 1.7200 6.3850 1.7200 6.3850 1.6900 5.5750 1.6900 5.5750 1.5700 6.3850 1.5700
                 6.3850 1.4800 6.5050 1.4800 ;
        POLYGON  6.1550 1.1200 5.9150 1.1200 5.9150 0.8500 5.2150 0.8500 5.2150 1.6900 4.7350 1.6900
                 4.7350 1.5700 5.0950 1.5700 5.0950 0.8500 4.7550 0.8500 4.7550 0.6800 4.9950 0.6800
                 4.9950 0.7300 6.0350 0.7300 6.0350 1.0000 6.1550 1.0000 ;
        RECT  3.1450 2.0500 5.6550 2.1700 ;
        POLYGON  4.3750 1.6900 4.1350 1.6900 4.1350 1.5700 4.1550 1.5700 4.1550 0.8500 2.8950 0.8500
                 2.8950 0.4800 2.7350 0.4800 2.7350 0.3600 3.0150 0.3600 3.0150 0.7300 4.1550 0.7300
                 4.1550 0.6200 4.2750 0.6200 4.2750 1.5700 4.3750 1.5700 ;
        POLYGON  3.7550 1.1400 3.4550 1.1400 3.4550 1.1100 2.7950 1.1100 2.7950 1.5700 3.2250 1.5700
                 3.2250 1.6900 2.6750 1.6900 2.6750 1.1100 2.6550 1.1100 2.6550 0.7400 2.4950 0.7400
                 2.4950 0.5600 2.1350 0.5600 2.1350 1.2000 1.5750 1.2000 1.5750 1.0800 2.0150 1.0800
                 2.0150 0.4400 2.6150 0.4400 2.6150 0.6200 2.7750 0.6200 2.7750 0.9900 3.5750 0.9900
                 3.5750 1.0200 3.7550 1.0200 ;
        POLYGON  1.2150 1.5800 1.0950 1.5800 1.0950 1.4600 0.9850 1.4600 0.9850 1.1800 0.3750 1.1800
                 0.3750 1.0600 0.9850 1.0600 0.9850 0.6800 1.1050 0.6800 1.1050 1.3400 1.2150 1.3400 ;
    END
END SDFFRXL

MACRO SDFFRX4
    CLASS CORE ;
    FOREIGN SDFFRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.6300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6150 0.3600 1.7350 1.5300 ;
        RECT  0.8950 0.3600 1.7350 0.4800 ;
        RECT  0.9200 0.9200 1.2350 1.0400 ;
        RECT  0.3900 0.9000 1.0400 1.0200 ;
        RECT  0.8950 0.3600 1.0150 1.0200 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        RECT  0.3900 0.9000 0.5100 1.4350 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1600 0.8350 1.5300 ;
        RECT  0.6500 1.1400 0.8000 1.5300 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9350 1.2900 2.2500 1.4350 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.9350 1.2900 2.0550 1.5300 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0600 2.5400 1.5300 ;
        RECT  2.3700 0.9600 2.4900 1.4600 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8350 1.0000 8.9550 1.2400 ;
        RECT  7.7950 1.0000 8.9550 1.1200 ;
        RECT  7.9150 0.5700 8.0350 1.1200 ;
        RECT  7.1950 0.5700 8.0350 0.6900 ;
        RECT  7.1950 0.3800 7.3150 0.6900 ;
        RECT  6.2950 0.3800 7.3150 0.5000 ;
        RECT  5.3850 1.2400 6.4150 1.3600 ;
        RECT  6.2950 0.3800 6.4150 1.3600 ;
        RECT  6.2450 0.9400 6.4150 1.3600 ;
        RECT  6.1050 0.9400 6.4150 1.0900 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7150 1.4400 10.8350 2.2100 ;
        RECT  10.5350 1.4400 10.8350 1.5600 ;
        RECT  9.4750 0.6800 10.6750 0.8000 ;
        RECT  9.9300 1.3200 10.6550 1.4400 ;
        RECT  9.9300 1.1750 10.0800 1.4400 ;
        RECT  9.9300 0.6800 10.0500 1.5600 ;
        RECT  9.8750 1.4400 9.9950 2.2100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.3950 0.6800 12.5950 0.8000 ;
        RECT  12.3950 1.4400 12.5150 2.2100 ;
        RECT  12.2150 1.4400 12.5150 1.5600 ;
        RECT  11.6700 1.3200 12.3350 1.4400 ;
        RECT  11.6700 1.1750 11.8200 1.4400 ;
        RECT  11.6700 0.6800 11.7900 1.5600 ;
        RECT  11.5550 1.4400 11.6750 2.2100 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.6300 0.1800 ;
        RECT  12.8350 -0.1800 13.0750 0.3200 ;
        RECT  11.8750 -0.1800 12.1150 0.3200 ;
        RECT  10.9150 -0.1800 11.1550 0.3200 ;
        RECT  9.9550 -0.1800 10.1950 0.3200 ;
        RECT  8.9950 -0.1800 9.2350 0.3200 ;
        RECT  7.5950 0.3300 7.8350 0.4500 ;
        RECT  7.5950 -0.1800 7.7150 0.4500 ;
        RECT  5.8750 0.6800 6.1750 0.8000 ;
        RECT  6.0550 -0.1800 6.1750 0.8000 ;
        RECT  2.9550 -0.1800 3.0750 0.9200 ;
        RECT  1.8950 -0.1800 2.0150 0.7800 ;
        RECT  0.5550 -0.1800 0.6750 0.7800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.6300 2.7900 ;
        RECT  12.8150 1.5600 12.9350 2.7900 ;
        RECT  11.9750 1.5600 12.0950 2.7900 ;
        RECT  11.1350 1.5600 11.2550 2.7900 ;
        RECT  10.2950 1.5600 10.4150 2.7900 ;
        RECT  9.4550 1.5600 9.5750 2.7900 ;
        RECT  8.3150 1.7200 8.4350 2.7900 ;
        RECT  7.4150 1.7200 7.6550 2.0900 ;
        RECT  7.4150 1.7200 7.5350 2.7900 ;
        RECT  5.9350 2.1700 6.0550 2.7900 ;
        RECT  5.8150 2.1700 6.0550 2.2900 ;
        RECT  4.7350 2.2000 4.9750 2.7900 ;
        RECT  3.1400 2.0000 3.2600 2.7900 ;
        RECT  2.0950 1.8900 2.2150 2.7900 ;
        RECT  0.6350 1.8900 0.7550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.4950 0.8600 13.3550 0.8600 13.3550 2.2100 13.2350 2.2100 13.2350 1.4400
                 12.6550 1.4400 12.6550 1.2000 12.7750 1.2000 12.7750 1.3200 13.2350 1.3200
                 13.2350 0.7400 13.3750 0.7400 13.3750 0.6200 13.4950 0.6200 ;
        POLYGON  13.0950 1.2000 12.9750 1.2000 12.9750 0.5600 10.9150 0.5600 10.9150 1.0600
                 10.8950 1.0600 10.8950 1.1800 10.7750 1.1800 10.7750 0.9400 10.7950 0.9400
                 10.7950 0.5600 8.4750 0.5600 8.4750 0.7600 8.3550 0.7600 8.3550 0.4400 13.0950 0.4400 ;
        POLYGON  9.3350 1.6000 8.8550 1.6000 8.8550 2.1500 8.7350 2.1500 8.7350 1.6000 8.0150 1.6000
                 8.0150 2.1500 7.8950 2.1500 7.8950 1.6000 7.3150 1.6000 7.3150 1.3100 7.4350 1.3100
                 7.4350 1.4800 9.2150 1.4800 9.2150 1.2200 9.3350 1.2200 ;
        POLYGON  8.3750 1.3600 7.5550 1.3600 7.5550 0.9300 6.9150 0.9300 6.9150 1.8100 6.9550 1.8100
                 6.9550 1.9300 6.7150 1.9300 6.7150 1.8100 6.7950 1.8100 6.7950 0.7400 6.9550 0.7400
                 6.9550 0.6200 7.0750 0.6200 7.0750 0.8100 7.6750 0.8100 7.6750 1.2400 8.3750 1.2400 ;
        POLYGON  7.2750 1.1700 7.1950 1.1700 7.1950 2.1700 6.8150 2.1700 6.8150 2.2500 6.5750 2.2500
                 6.5750 2.1700 6.1750 2.1700 6.1750 2.0500 5.6950 2.0500 5.6950 2.2000 5.0950 2.2000
                 5.0950 2.0800 4.3450 2.0800 4.3450 2.0600 4.3350 2.0600 4.3350 2.0000 3.4200 2.0000
                 3.4200 1.8800 4.3450 1.8800 4.3450 1.8200 4.4650 1.8200 4.4650 1.9600 5.2150 1.9600
                 5.2150 2.0800 5.5750 2.0800 5.5750 1.9300 6.2950 1.9300 6.2950 2.0500 7.0750 2.0500
                 7.0750 1.1700 7.0350 1.1700 7.0350 1.0500 7.2750 1.0500 ;
        POLYGON  6.6550 1.6900 6.5350 1.6900 6.5350 1.8100 6.2950 1.8100 6.2950 1.6000 5.0850 1.6000
                 5.0850 1.3100 5.2050 1.3100 5.2050 1.4800 6.5350 1.4800 6.5350 0.6200 6.6550 0.6200 ;
        POLYGON  5.9850 1.1200 4.8450 1.1200 4.8450 1.2200 4.4850 1.2200 4.4850 1.5800 4.3050 1.5800
                 4.3050 1.7000 4.1850 1.7000 4.1850 1.4600 4.3650 1.4600 4.3650 1.1000 4.7250 1.1000
                 4.7250 0.6200 4.8450 0.6200 4.8450 1.0000 5.9850 1.0000 ;
        POLYGON  5.9350 0.4800 4.4150 0.4800 4.4150 0.5000 4.1500 0.5000 4.1500 0.7400 3.8850 0.7400
                 3.8850 0.9800 4.0050 0.9800 4.0050 1.1000 3.7650 1.1000 3.7650 0.9800 3.5550 0.9800
                 3.5550 1.5200 3.3150 1.5200 3.3150 1.4000 3.4350 1.4000 3.4350 0.8600 3.3150 0.8600
                 3.3150 0.7400 3.5550 0.7400 3.5550 0.8600 3.7650 0.8600 3.7650 0.6200 4.0300 0.6200
                 4.0300 0.3800 4.2950 0.3800 4.2950 0.3600 5.9350 0.3600 ;
        POLYGON  5.4550 1.9600 5.3350 1.9600 5.3350 1.8400 4.6050 1.8400 4.6050 1.3400 4.7250 1.3400
                 4.7250 1.7200 5.4550 1.7200 ;
        POLYGON  4.4250 0.9800 4.2450 0.9800 4.2450 1.3400 3.8850 1.3400 3.8850 1.7600 3.0200 1.7600
                 3.0200 2.2500 2.3350 2.2500 2.3350 1.7700 1.8000 1.7700 1.8000 1.8900 1.5350 1.8900
                 1.5350 2.0100 1.4150 2.0100 1.4150 1.8900 1.3750 1.8900 1.3750 0.7200 1.1350 0.7200
                 1.1350 0.6000 1.4950 0.6000 1.4950 1.7700 1.6800 1.7700 1.6800 1.6500 2.4550 1.6500
                 2.4550 2.1300 2.9000 2.1300 2.9000 1.6400 3.7650 1.6400 3.7650 1.2200 4.1250 1.2200
                 4.1250 0.8600 4.3050 0.8600 4.3050 0.6200 4.4250 0.6200 ;
        POLYGON  3.2750 1.2000 2.7800 1.2000 2.7800 1.7700 2.6950 1.7700 2.6950 2.0100 2.5750 2.0100
                 2.5750 1.6500 2.6600 1.6500 2.6600 0.8400 2.3150 0.8400 2.3150 0.5400 2.4350 0.5400
                 2.4350 0.7200 2.7800 0.7200 2.7800 1.0800 3.2750 1.0800 ;
        POLYGON  1.2550 1.7700 0.3350 1.7700 0.3350 2.0100 0.2150 2.0100 0.2150 1.8900 0.1200 1.8900
                 0.1200 0.9350 0.1350 0.9350 0.1350 0.5400 0.2550 0.5400 0.2550 1.0550 0.2400 1.0550
                 0.2400 1.6500 1.1350 1.6500 1.1350 1.4500 1.2550 1.4500 ;
    END
END SDFFRX4

MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.8700 2.8850 1.1000 ;
        RECT  2.6950 0.8700 2.8150 1.2800 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7600 2.0500 6.3250 2.1700 ;
        RECT  4.7600 1.8700 4.8800 2.1700 ;
        RECT  4.6850 1.4350 4.8050 1.9900 ;
        RECT  4.1300 1.4350 4.8050 1.5550 ;
        RECT  4.1300 1.1750 4.2800 1.5550 ;
        RECT  3.9450 1.1700 4.2500 1.2900 ;
        END
    END RN
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7700 1.1750 9.0850 1.3200 ;
        RECT  8.9650 1.0800 9.0850 1.3200 ;
        RECT  8.7700 1.1750 8.9200 1.4350 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.0250 1.3000 10.3050 1.4200 ;
        RECT  9.8750 1.8100 10.1450 1.9600 ;
        RECT  10.0250 1.3000 10.1450 1.9600 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5100 1.1750 10.6600 1.4350 ;
        RECT  9.7850 1.0600 10.6300 1.1800 ;
        RECT  10.5100 1.0550 10.6300 1.4350 ;
        RECT  9.7850 1.0600 9.9050 1.5000 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1950 0.8850 1.3800 1.1450 ;
        RECT  1.0350 1.4000 1.3150 1.5200 ;
        RECT  1.1950 0.5900 1.3150 1.5200 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0350 0.8850 2.2500 1.1450 ;
        RECT  1.9950 1.4000 2.2350 1.5200 ;
        RECT  2.0350 0.5900 2.1550 1.5200 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.2250 -0.1800 10.4650 0.3800 ;
        RECT  8.8250 -0.1800 8.9450 0.9200 ;
        RECT  5.9250 -0.1800 6.1650 0.3200 ;
        RECT  4.0650 0.4500 4.3050 0.5700 ;
        RECT  4.1850 -0.1800 4.3050 0.5700 ;
        RECT  2.4550 -0.1800 2.5750 0.6400 ;
        RECT  1.6150 -0.1800 1.7350 0.6400 ;
        RECT  0.7750 -0.1800 0.8950 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.2850 2.2200 10.4050 2.7900 ;
        RECT  8.8850 2.2200 9.0050 2.7900 ;
        RECT  6.7250 2.0500 6.9650 2.1700 ;
        RECT  6.7250 2.0500 6.8450 2.7900 ;
        RECT  5.7650 2.2900 6.0050 2.7900 ;
        RECT  4.1250 2.2300 4.2450 2.7900 ;
        RECT  3.2450 1.8800 3.3650 2.7900 ;
        RECT  2.5350 1.9800 2.6550 2.7900 ;
        RECT  1.5150 1.8800 1.7550 2.0000 ;
        RECT  1.5150 1.8800 1.6350 2.7900 ;
        RECT  0.5550 1.8800 0.7950 2.0000 ;
        RECT  0.5550 1.8800 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.9000 1.7000 10.8850 1.7000 10.8850 1.8200 10.7650 1.8200 10.7650 1.5800
                 10.7800 1.5800 10.7800 0.9200 10.7650 0.9200 10.7650 0.6800 10.3150 0.6800
                 10.3150 0.6200 9.4050 0.6200 9.4050 1.2400 9.4250 1.2400 9.4250 1.4800 9.2850 1.4800
                 9.2850 0.5000 9.6650 0.5000 9.6650 0.4200 9.9050 0.4200 9.9050 0.5000 10.4350 0.5000
                 10.4350 0.5600 10.8850 0.5600 10.8850 0.8000 10.9000 0.8000 ;
        POLYGON  9.7650 0.8600 9.6650 0.8600 9.6650 1.7600 9.6250 1.7600 9.6250 2.0000 8.1050 2.0000
                 8.1050 1.7000 8.0150 1.7000 8.0150 1.3400 7.7150 1.3400 7.7150 0.8600 7.4250 0.8600
                 7.4250 0.6200 7.5450 0.6200 7.5450 0.7400 7.8350 0.7400 7.8350 1.2200 8.1350 1.2200
                 8.1350 1.5800 8.2250 1.5800 8.2250 1.8800 9.5050 1.8800 9.5050 1.6400 9.5450 1.6400
                 9.5450 0.8600 9.5250 0.8600 9.5250 0.7400 9.7650 0.7400 ;
        POLYGON  8.7450 2.2400 7.8650 2.2400 7.8650 1.9400 7.4550 1.9400 7.4550 2.0400 7.3350 2.0400
                 7.3350 1.9400 7.2850 1.9400 7.2850 1.9300 5.1650 1.9300 5.1650 1.0750 5.1250 1.0750
                 5.1250 0.5600 4.5800 0.5600 4.5800 0.8100 3.6650 0.8100 3.6650 0.5000 3.0550 0.5000
                 3.0550 0.6300 3.1250 0.6300 3.1250 1.5200 2.8750 1.5200 2.8750 1.4000 3.0050 1.4000
                 3.0050 0.7500 2.9350 0.7500 2.9350 0.3800 3.7850 0.3800 3.7850 0.6900 4.4600 0.6900
                 4.4600 0.4400 4.6250 0.4400 4.6250 0.3600 4.8650 0.3600 4.8650 0.4400 5.2450 0.4400
                 5.2450 0.9550 5.2850 0.9550 5.2850 1.8100 7.3350 1.8100 7.3350 1.8000 7.4550 1.8000
                 7.4550 1.8200 7.9850 1.8200 7.9850 2.1200 8.7450 2.1200 ;
        POLYGON  8.5850 1.7600 8.3450 1.7600 8.3450 1.6400 8.4050 1.6400 8.4050 0.9800 8.0750 0.9800
                 8.0750 1.1000 7.9550 1.1000 7.9550 0.5000 6.4050 0.5000 6.4050 0.5600 5.4850 0.5600
                 5.4850 0.4800 5.3650 0.4800 5.3650 0.3600 5.6050 0.3600 5.6050 0.4400 6.2850 0.4400
                 6.2850 0.3800 6.8050 0.3800 6.8050 0.3600 7.0450 0.3600 7.0450 0.3800 8.0750 0.3800
                 8.0750 0.8600 8.4050 0.8600 8.4050 0.6800 8.5250 0.6800 8.5250 1.6400 8.5850 1.6400 ;
        POLYGON  7.7150 1.7000 7.5950 1.7000 7.5950 1.5800 7.4750 1.5800 7.4750 1.3800 5.8450 1.3800
                 5.8450 1.3700 5.7250 1.3700 5.7250 1.2500 5.9650 1.2500 5.9650 1.2600 7.0050 1.2600
                 7.0050 0.6200 7.1250 0.6200 7.1250 1.2600 7.5950 1.2600 7.5950 1.4600 7.7150 1.4600 ;
        POLYGON  7.3550 1.6400 6.4850 1.6400 6.4850 1.6900 6.2450 1.6900 6.2450 1.5700 6.3650 1.5700
                 6.3650 1.5200 7.3550 1.5200 ;
        POLYGON  6.7050 1.1400 6.4650 1.1400 6.4650 1.1300 5.6050 1.1300 5.6050 1.5700 5.6450 1.5700
                 5.6450 1.6900 5.4050 1.6900 5.4050 1.5700 5.4850 1.5700 5.4850 0.8000 5.3650 0.8000
                 5.3650 0.6800 5.6050 0.6800 5.6050 1.0100 6.5850 1.0100 6.5850 1.0200 6.7050 1.0200 ;
        POLYGON  5.0450 1.7500 4.9250 1.7500 4.9250 1.3150 4.7650 1.3150 4.7650 1.0500 3.8250 1.0500
                 3.8250 1.1400 3.5250 1.1400 3.5250 1.0200 3.7050 1.0200 3.7050 0.9300 4.7650 0.9300
                 4.7650 0.6800 5.0050 0.6800 5.0050 0.8000 4.8850 0.8000 4.8850 1.1950 5.0450 1.1950 ;
        POLYGON  4.5650 2.2100 4.4450 2.2100 4.4450 2.0700 3.7250 2.0700 3.7250 1.5300 3.4050 1.5300
                 3.4050 1.7600 0.5550 1.7600 0.5550 1.0000 0.6750 1.0000 0.6750 1.6400 1.7550 1.6400
                 1.7550 1.0200 1.8750 1.0200 1.8750 1.6400 2.3700 1.6400 2.3700 1.0000 2.4900 1.0000
                 2.4900 1.6400 3.2850 1.6400 3.2850 0.7800 3.4250 0.7800 3.4250 0.6200 3.5450 0.6200
                 3.5450 0.9000 3.4050 0.9000 3.4050 1.4100 3.8450 1.4100 3.8450 1.9500 4.5650 1.9500 ;
        POLYGON  1.0550 1.1700 0.9350 1.1700 0.9350 0.8800 0.4150 0.8800 0.4150 1.4600 0.2550 1.4600
                 0.2550 1.5800 0.1350 1.5800 0.1350 1.3400 0.2950 1.3400 0.2950 0.5900 0.4150 0.5900
                 0.4150 0.7600 1.0550 0.7600 ;
    END
END SDFFRX2

MACRO SDFFRX1
    CLASS CORE ;
    FOREIGN SDFFRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.7300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8450 1.3400 2.1250 1.4600 ;
        RECT  2.0050 1.2200 2.1250 1.4600 ;
        RECT  1.8100 1.4650 1.9650 1.7250 ;
        RECT  1.8450 1.3400 1.9650 1.7250 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3456  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 2.8800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2050 1.2050 3.5250 1.4250 ;
        RECT  3.2050 1.2050 3.4650 1.4500 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1900 0.7600 8.4450 0.9600 ;
        RECT  8.1900 0.7600 8.3400 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5850 0.9400 9.8450 1.1700 ;
        RECT  9.6650 0.9400 9.7850 1.3500 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.0050 0.8850 10.3700 1.1450 ;
        RECT  10.0050 0.7000 10.1250 1.1450 ;
        RECT  9.3450 0.7000 10.1250 0.8200 ;
        RECT  8.8050 1.0300 9.4650 1.1500 ;
        RECT  9.3450 0.7000 9.4650 1.1500 ;
        RECT  8.8050 1.0300 8.9250 1.2700 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 2.2100 ;
        RECT  1.2300 0.8850 1.4850 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.7300 0.1800 ;
        RECT  9.7650 0.4600 10.0050 0.5800 ;
        RECT  9.7650 -0.1800 9.8850 0.5800 ;
        RECT  8.3250 -0.1800 8.4450 0.6400 ;
        RECT  5.7650 0.4700 6.0050 0.5900 ;
        RECT  5.8850 -0.1800 6.0050 0.5900 ;
        RECT  3.5450 -0.1800 3.6650 0.6050 ;
        RECT  1.7250 0.5500 1.9650 0.6700 ;
        RECT  1.7250 -0.1800 1.8450 0.6700 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.7300 2.7900 ;
        RECT  9.7250 1.7100 9.8450 2.7900 ;
        RECT  8.4850 2.2300 8.6050 2.7900 ;
        RECT  6.4450 2.0500 6.6850 2.1700 ;
        RECT  6.4450 2.0500 6.5650 2.7900 ;
        RECT  5.4850 2.2900 5.7250 2.7900 ;
        RECT  3.4850 2.2900 3.7250 2.7900 ;
        RECT  2.6550 2.1500 2.7750 2.7900 ;
        RECT  1.7850 1.8450 1.9050 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.6100 1.7100 10.2650 1.7100 10.2650 1.8300 10.1450 1.8300 10.1450 1.5900
                 9.2850 1.5900 9.2850 1.4500 9.1650 1.4500 9.1650 1.3300 9.4050 1.3300 9.4050 1.4700
                 10.4900 1.4700 10.4900 0.7650 10.2450 0.7650 10.2450 0.4000 10.3650 0.4000
                 10.3650 0.6450 10.6100 0.6450 ;
        POLYGON  9.3650 0.5800 9.2250 0.5800 9.2250 0.9100 8.6850 0.9100 8.6850 1.7700 9.2450 1.7700
                 9.2450 1.8900 8.6850 1.8900 8.6850 2.0100 7.6150 2.0100 7.6150 1.3400 7.4050 1.3400
                 7.4050 0.8600 7.3050 0.8600 7.3050 0.6200 7.4250 0.6200 7.4250 0.7400 7.5250 0.7400
                 7.5250 1.2200 7.7350 1.2200 7.7350 1.8900 8.5650 1.8900 8.5650 0.7900 9.1050 0.7900
                 9.1050 0.4600 9.3650 0.4600 ;
        POLYGON  8.3450 2.2500 7.2200 2.2500 7.2200 1.9400 7.0750 1.9400 7.0750 2.0400 6.9550 2.0400
                 6.9550 1.9300 2.2650 1.9300 2.2650 1.5700 2.3250 1.5700 2.3250 0.7400 2.5650 0.7400
                 2.5650 0.8600 2.4450 0.8600 2.4450 1.6900 2.3850 1.6900 2.3850 1.8100 4.1050 1.8100
                 4.1050 0.9400 4.2250 0.9400 4.2250 1.8100 4.7650 1.8100 4.7650 1.3700 4.6250 1.3700
                 4.6250 1.2500 4.8850 1.2500 4.8850 1.8100 6.9550 1.8100 6.9550 1.8000 7.0750 1.8000
                 7.0750 1.8200 7.3400 1.8200 7.3400 2.1300 8.3450 2.1300 ;
        POLYGON  8.1850 1.7700 7.9450 1.7700 7.9450 0.9800 7.7650 0.9800 7.7650 1.1000 7.6450 1.1000
                 7.6450 0.5000 6.2450 0.5000 6.2450 0.8300 5.5250 0.8300 5.5250 0.5000 5.1650 0.5000
                 5.1650 1.1800 5.0450 1.1800 5.0450 0.3800 5.6450 0.3800 5.6450 0.7100 6.1250 0.7100
                 6.1250 0.3800 6.5450 0.3800 6.5450 0.3600 6.7850 0.3600 6.7850 0.3800 7.7650 0.3800
                 7.7650 0.4000 7.8850 0.4000 7.8850 0.8600 8.0650 0.8600 8.0650 1.6500 8.1850 1.6500 ;
        POLYGON  7.3150 1.7000 7.1950 1.7000 7.1950 1.5800 7.1650 1.5800 7.1650 1.4000 5.6450 1.4000
                 5.6450 1.4300 5.5250 1.4300 5.5250 1.1900 5.6450 1.1900 5.6450 1.2800 6.8850 1.2800
                 6.8850 0.6200 7.0050 0.6200 7.0050 1.2800 7.2850 1.2800 7.2850 1.4600 7.3150 1.4600 ;
        POLYGON  6.9550 1.6400 6.2050 1.6400 6.2050 1.6900 5.9650 1.6900 5.9650 1.5700 6.0850 1.5700
                 6.0850 1.5200 6.9550 1.5200 ;
        POLYGON  6.5650 1.1200 6.3250 1.1200 6.3250 1.0700 5.4050 1.0700 5.4050 1.6900 5.0050 1.6900
                 5.0050 1.5700 5.2850 1.5700 5.2850 0.6200 5.4050 0.6200 5.4050 0.9500 6.4450 0.9500
                 6.4450 1.0000 6.5650 1.0000 ;
        RECT  3.1650 2.0500 6.0450 2.1700 ;
        POLYGON  4.6450 1.6900 4.3850 1.6900 4.3850 0.8200 3.9750 0.8200 3.9750 0.8450 3.0850 0.8450
                 3.0850 0.4800 2.9250 0.4800 2.9250 0.3600 3.2050 0.3600 3.2050 0.7250 3.8550 0.7250
                 3.8550 0.7000 4.3850 0.7000 4.3850 0.6200 4.5050 0.6200 4.5050 1.5700 4.6450 1.5700 ;
        POLYGON  3.8850 1.2050 3.7650 1.2050 3.7650 1.0850 3.0850 1.0850 3.0850 1.5700 3.2450 1.5700
                 3.2450 1.6900 2.9650 1.6900 2.9650 1.0850 2.8450 1.0850 2.8450 0.7400 2.6850 0.7400
                 2.6850 0.6200 2.2050 0.6200 2.2050 1.1000 1.7250 1.1000 1.7250 1.2400 1.6050 1.2400
                 1.6050 0.9800 2.0850 0.9800 2.0850 0.5000 2.8050 0.5000 2.8050 0.6200 2.9650 0.6200
                 2.9650 0.9650 3.8850 0.9650 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END SDFFRX1

MACRO SDFFRHQX8
    CLASS CORE ;
    FOREIGN SDFFRHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.9200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7750 0.6650 2.8950 0.9600 ;
        RECT  2.6550 0.8400 2.7750 2.0850 ;
        RECT  0.2550 1.0250 2.7750 1.1450 ;
        RECT  1.9350 0.6650 2.0550 1.1450 ;
        RECT  1.8150 0.9050 1.9350 2.0850 ;
        RECT  1.0950 0.6650 1.2150 1.1450 ;
        RECT  0.9750 0.9050 1.0950 2.0800 ;
        RECT  0.2550 0.8850 0.5100 1.1450 ;
        RECT  0.2550 0.6650 0.3750 1.2650 ;
        RECT  0.1350 1.1450 0.2550 2.0800 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.4020  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4100  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.9805  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4150 0.9800 4.6950 1.1000 ;
        RECT  4.4150 0.3600 4.5350 1.1000 ;
        RECT  3.6350 0.3600 4.5350 0.4800 ;
        RECT  3.3750 1.0000 3.7550 1.1200 ;
        RECT  3.6350 0.3600 3.7550 1.1200 ;
        RECT  3.4950 0.9400 3.7550 1.1200 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1050 1.1850 6.3650 1.4100 ;
        RECT  6.2450 1.0100 6.3650 1.4100 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.5250 0.9300 11.6450 1.1700 ;
        RECT  11.0900 0.9300 11.6450 1.0500 ;
        RECT  11.0900 0.8850 11.2400 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.7400 1.2300 13.0550 1.4300 ;
        RECT  12.7400 1.2100 13.0350 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.1550 0.9900 13.3950 1.1100 ;
        RECT  12.0050 0.9700 13.3250 1.0900 ;
        RECT  13.0650 0.9400 13.3250 1.0900 ;
        RECT  12.0050 0.9700 12.1250 1.4400 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.9200 0.1800 ;
        RECT  13.0650 -0.1800 13.1850 0.8200 ;
        RECT  11.5250 -0.1800 11.6450 0.6400 ;
        RECT  8.5850 0.4300 8.8250 0.5500 ;
        RECT  8.7050 -0.1800 8.8250 0.5500 ;
        RECT  6.3250 -0.1800 6.5650 0.4100 ;
        RECT  4.7550 -0.1800 4.8750 0.6500 ;
        RECT  3.1950 -0.1800 3.3150 0.6500 ;
        RECT  2.3550 -0.1800 2.4750 0.6550 ;
        RECT  1.5150 -0.1800 1.6350 0.6550 ;
        RECT  0.6750 -0.1800 0.7950 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.9200 2.7900 ;
        RECT  12.9050 1.7950 13.0250 2.7900 ;
        RECT  11.4050 2.2800 11.6450 2.7900 ;
        RECT  9.3050 2.2600 9.5450 2.7900 ;
        RECT  8.4050 1.7500 8.5250 2.7900 ;
        RECT  6.3850 2.2500 6.6250 2.7900 ;
        RECT  5.5950 2.2500 5.8350 2.7900 ;
        RECT  4.7550 1.7000 4.8750 1.9900 ;
        RECT  4.7350 1.8700 4.8550 2.7900 ;
        RECT  3.9150 1.7000 4.0350 2.7900 ;
        RECT  3.0750 1.7000 3.1950 2.7900 ;
        RECT  2.2350 1.3400 2.3550 2.7900 ;
        RECT  1.3950 1.3400 1.5150 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.6350 1.6800 13.5050 1.6800 13.5050 1.8000 13.3850 1.8000 13.3850 1.6750
                 12.4050 1.6750 12.4050 1.2400 12.5250 1.2400 12.5250 1.5550 13.5150 1.5550
                 13.5150 0.8200 13.4850 0.8200 13.4850 0.5800 13.6050 0.5800 13.6050 0.7000
                 13.6350 0.7000 ;
        POLYGON  12.5450 0.8500 11.8850 0.8500 11.8850 1.5600 12.2850 1.5600 12.2850 2.2100
                 12.1650 2.2100 12.1650 1.6800 11.8850 1.6800 11.8850 1.8000 11.6200 1.8000
                 11.6200 1.9800 10.5950 1.9800 10.5950 1.3000 10.1350 1.3000 10.1350 0.7200
                 10.0850 0.7200 10.0850 0.6000 10.3250 0.6000 10.3250 0.7200 10.2550 0.7200
                 10.2550 1.1800 10.7150 1.1800 10.7150 1.8600 11.5000 1.8600 11.5000 1.6800
                 11.7650 1.6800 11.7650 0.7300 12.4250 0.7300 12.4250 0.5900 12.5450 0.5900 ;
        POLYGON  11.2850 2.2200 9.7200 2.2200 9.7200 2.1400 8.6450 2.1400 8.6450 1.6300 8.2850 1.6300
                 8.2850 2.0100 6.9850 2.0100 6.9850 1.8900 6.9250 1.8900 6.9250 0.8900 5.9650 0.8900
                 5.9650 1.5300 6.2250 1.5300 6.2250 1.6500 5.8450 1.6500 5.8450 0.7200 5.7250 0.7200
                 5.7250 0.6000 5.9650 0.6000 5.9650 0.7700 7.0450 0.7700 7.0450 1.7700 7.1050 1.7700
                 7.1050 1.8900 7.4650 1.8900 7.4650 1.1300 7.5850 1.1300 7.5850 1.8900 8.1650 1.8900
                 8.1650 1.5100 8.7650 1.5100 8.7650 2.0200 9.8400 2.0200 9.8400 2.1000 11.2850 2.1000 ;
        POLYGON  11.1650 1.7400 10.8500 1.7400 10.8500 1.0600 10.3750 1.0600 10.3750 0.9400
                 10.4950 0.9400 10.4950 0.4800 9.5450 0.4800 9.5450 0.8600 9.6450 0.8600 9.6450 1.1000
                 9.4250 1.1000 9.4250 0.7900 8.3450 0.7900 8.3450 0.4800 7.8650 0.4800 7.8650 0.9200
                 7.9850 0.9200 7.9850 1.0400 7.7450 1.0400 7.7450 0.3600 8.4650 0.3600 8.4650 0.6700
                 9.4250 0.6700 9.4250 0.3600 10.6150 0.3600 10.6150 0.9400 10.8500 0.9400
                 10.8500 0.5900 10.9700 0.5900 10.9700 1.6200 11.1650 1.6200 ;
        POLYGON  10.2950 1.9400 10.1750 1.9400 10.1750 1.5400 9.7650 1.5400 9.7650 1.3900 8.4650 1.3900
                 8.4650 1.3100 8.3450 1.3100 8.3450 1.1900 8.5850 1.1900 8.5850 1.2700 9.7650 1.2700
                 9.7650 0.7200 9.6650 0.7200 9.6650 0.6000 9.9050 0.6000 9.9050 0.7200 9.8850 0.7200
                 9.8850 1.4200 10.2950 1.4200 ;
        POLYGON  9.8750 1.9000 8.8850 1.9000 8.8850 1.5100 9.0050 1.5100 9.0050 1.7800 9.7550 1.7800
                 9.7550 1.6600 9.8750 1.6600 ;
        POLYGON  9.3050 1.1500 9.1850 1.1500 9.1850 1.0700 8.2250 1.0700 8.2250 1.2800 8.0450 1.2800
                 8.0450 1.7700 7.9250 1.7700 7.9250 1.1600 8.1050 1.1600 8.1050 0.7200 7.9850 0.7200
                 7.9850 0.6000 8.2250 0.6000 8.2250 0.9500 9.1850 0.9500 9.1850 0.9100 9.3050 0.9100 ;
        POLYGON  8.0850 2.2500 6.7450 2.2500 6.7450 2.1300 5.2150 2.1300 5.2150 2.2500 4.9750 2.2500
                 4.9750 2.1300 5.0950 2.1300 5.0950 2.0100 6.8650 2.0100 6.8650 2.1300 8.0850 2.1300 ;
        POLYGON  7.3450 1.7700 7.2250 1.7700 7.2250 0.6500 6.0850 0.6500 6.0850 0.4800 5.4800 0.4800
                 5.4800 0.5400 5.2150 0.5400 5.2150 1.0800 5.4350 1.0800 5.4350 1.2000 5.2150 1.2000
                 5.2150 1.3400 4.1750 1.3400 4.1750 1.0000 4.2950 1.0000 4.2950 1.2200 5.0950 1.2200
                 5.0950 0.4200 5.3600 0.4200 5.3600 0.3600 6.2050 0.3600 6.2050 0.5300 7.3450 0.5300 ;
        POLYGON  6.7250 1.8900 5.5550 1.8900 5.5550 1.5800 5.2950 1.5800 5.2950 1.8900 5.1750 1.8900
                 5.1750 1.5800 4.4550 1.5800 4.4550 1.9900 4.3350 1.9900 4.3350 1.5800 3.6150 1.5800
                 3.6150 1.9900 3.4950 1.9900 3.4950 1.5800 3.0150 1.5800 3.0150 1.2000 2.8950 1.2000
                 2.8950 1.0800 3.1350 1.0800 3.1350 1.4600 3.4950 1.4600 3.4950 1.3400 3.6150 1.3400
                 3.6150 1.4600 3.9150 1.4600 3.9150 0.6000 4.0350 0.6000 4.0350 1.4600 5.5550 1.4600
                 5.5550 0.9600 5.3350 0.9600 5.3350 0.6600 5.5750 0.6600 5.5750 0.8400 5.6750 0.8400
                 5.6750 1.7700 6.6050 1.7700 6.6050 1.1300 6.7250 1.1300 ;
    END
END SDFFRHQX8

MACRO SDFFRHQX4
    CLASS CORE ;
    FOREIGN SDFFRHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0800 0.6900 2.4400 0.8100 ;
        RECT  1.9950 1.4900 2.2350 1.6100 ;
        RECT  2.0800 0.6900 2.2000 1.6100 ;
        RECT  1.2300 0.8850 2.2000 1.0050 ;
        RECT  1.2600 0.7650 1.5400 1.0050 ;
        RECT  1.4200 0.6300 1.5400 1.0050 ;
        RECT  1.0350 1.4900 1.3800 1.6100 ;
        RECT  1.2600 0.7650 1.3800 1.6100 ;
        RECT  1.2300 0.8850 1.3800 1.1450 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.9800 0.5100 1.4350 ;
        RECT  0.3900 0.9300 0.5100 1.4350 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2580  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7150 1.0900 6.8350 1.3300 ;
        RECT  6.1350 1.2200 6.7350 1.3400 ;
        RECT  6.6150 1.2100 6.8350 1.3300 ;
        RECT  6.1350 0.3600 6.2550 1.3400 ;
        RECT  5.0550 0.3600 6.2550 0.4800 ;
        RECT  3.7350 0.4700 5.1750 0.5900 ;
        RECT  3.9350 0.4700 4.0550 1.1000 ;
        RECT  2.9400 0.3600 3.8550 0.4800 ;
        RECT  2.6800 0.8850 3.0600 1.1250 ;
        RECT  2.9400 0.3600 3.0600 1.1250 ;
        RECT  2.6800 0.8850 2.8300 1.1450 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.9050 0.9700 10.0250 1.2100 ;
        RECT  9.5850 0.9700 10.0250 1.0900 ;
        RECT  9.5850 0.9400 9.8450 1.0900 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0900 1.0200 11.2650 1.4400 ;
        RECT  11.1450 1.0000 11.2650 1.4400 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6150 1.2300 11.8750 1.3800 ;
        RECT  11.6150 1.0700 11.7650 1.3800 ;
        RECT  11.5250 0.7600 11.6450 1.1900 ;
        RECT  10.6050 0.7600 11.6450 0.8800 ;
        RECT  10.6050 0.7600 10.8450 1.0900 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.2850 -0.1800 11.4050 0.6400 ;
        RECT  9.6850 0.4600 9.9250 0.5800 ;
        RECT  9.6850 -0.1800 9.8050 0.5800 ;
        RECT  6.5550 -0.1800 6.6750 0.6800 ;
        RECT  4.3950 -0.1800 4.6350 0.3500 ;
        RECT  2.6800 -0.1800 2.8000 0.6800 ;
        RECT  1.8400 -0.1800 1.9600 0.6800 ;
        RECT  1.0000 -0.1800 1.1200 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.2850 1.8000 11.4050 2.7900 ;
        RECT  9.9850 1.8500 10.1050 2.7900 ;
        RECT  9.9700 1.6900 10.0900 1.9700 ;
        RECT  7.6750 2.2100 7.9150 2.7900 ;
        RECT  6.4350 2.2100 6.6750 2.7900 ;
        RECT  4.4550 2.2300 4.5750 2.7900 ;
        RECT  3.4950 2.2300 3.6150 2.7900 ;
        RECT  2.4750 1.9700 2.7150 2.0900 ;
        RECT  2.4750 1.9700 2.5950 2.7900 ;
        RECT  1.5150 1.9700 1.7550 2.0900 ;
        RECT  1.5150 1.9700 1.6350 2.7900 ;
        RECT  0.5550 1.9700 0.7950 2.0900 ;
        RECT  0.5550 1.9700 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.1150 1.7400 11.7050 1.7400 11.7050 1.6800 10.8500 1.6800 10.8500 1.4200
                 10.7250 1.4200 10.7250 1.3300 10.2250 1.3300 10.2250 0.9400 10.3450 0.9400
                 10.3450 1.2100 10.9650 1.2100 10.9650 1.3000 10.9700 1.3000 10.9700 1.5600
                 11.9950 1.5600 11.9950 0.9500 11.7650 0.9500 11.7650 0.5900 11.8850 0.5900
                 11.8850 0.8300 12.1150 0.8300 ;
        POLYGON  10.7300 2.2100 10.6100 2.2100 10.6100 1.6800 10.4850 1.6800 10.4850 1.5700
                 9.2750 1.5700 9.2750 1.5200 9.1550 1.5200 9.1550 1.4000 9.3450 1.4000 9.3450 0.5300
                 8.4350 0.5300 8.4350 0.6800 8.3150 0.6800 8.3150 0.4100 9.4650 0.4100 9.4650 0.7000
                 10.3250 0.7000 10.3250 0.5200 10.5650 0.5200 10.5650 0.6400 10.4450 0.6400
                 10.4450 0.8200 9.4650 0.8200 9.4650 1.4500 10.6050 1.4500 10.6050 1.5600
                 10.7300 1.5600 ;
        POLYGON  9.8650 2.2500 8.0750 2.2500 8.0750 2.0900 6.1500 2.0900 6.1500 2.1900 5.4750 2.1900
                 5.4750 2.2100 5.2350 2.2100 5.2350 2.1900 4.7050 2.1900 4.7050 2.1100 3.3150 2.1100
                 3.3150 1.8500 0.1350 1.8500 0.1350 1.6750 0.1200 1.6750 0.1200 0.6900 0.6350 0.6900
                 0.6350 0.8100 0.2400 0.8100 0.2400 1.5550 0.2550 1.5550 0.2550 1.7300 3.4350 1.7300
                 3.4350 1.9900 4.8250 1.9900 4.8250 2.0700 6.0300 2.0700 6.0300 1.9700 8.1950 1.9700
                 8.1950 2.1300 9.8650 2.1300 ;
        POLYGON  9.6450 1.9700 9.0350 1.9700 9.0350 2.0100 8.3150 2.0100 8.3150 1.8500 5.5350 1.8500
                 5.5350 1.3200 5.0150 1.3200 5.0150 1.0800 5.1350 1.0800 5.1350 1.2000 5.5350 1.2000
                 5.5350 0.9200 5.7750 0.9200 5.7750 1.0400 5.6550 1.0400 5.6550 1.7300 8.3150 1.7300
                 8.3150 1.1600 7.6950 1.1600 7.6950 1.0400 8.4350 1.0400 8.4350 1.8900 8.9150 1.8900
                 8.9150 0.6500 9.2250 0.6500 9.2250 0.7700 9.0350 0.7700 9.0350 1.8500 9.5250 1.8500
                 9.5250 1.7300 9.6450 1.7300 ;
        POLYGON  8.7950 1.7700 8.5550 1.7700 8.5550 0.9200 6.4950 0.9200 6.4950 1.1000 6.3750 1.1000
                 6.3750 0.8000 7.8950 0.8000 7.8950 0.5400 8.0150 0.5400 8.0150 0.8000 8.6750 0.8000
                 8.6750 1.4000 8.7950 1.4000 ;
        POLYGON  8.1950 1.6100 7.1950 1.6100 7.1950 1.4900 8.0750 1.4900 8.0750 1.3400 8.1950 1.3400 ;
        POLYGON  7.5750 1.2900 7.4550 1.2900 7.4550 1.3700 7.0750 1.3700 7.0750 1.5800 6.0150 1.5800
                 6.0150 1.6100 5.7750 1.6100 5.7750 1.4900 5.8950 1.4900 5.8950 0.7200 5.7750 0.7200
                 5.7750 0.6000 6.0150 0.6000 6.0150 1.4600 6.9550 1.4600 6.9550 1.2500 7.3350 1.2500
                 7.3350 1.1700 7.5750 1.1700 ;
        POLYGON  5.5950 0.7200 5.4150 0.7200 5.4150 0.8300 4.8950 0.8300 4.8950 1.4400 5.2750 1.4400
                 5.2750 1.9500 5.1550 1.9500 5.1550 1.5600 4.7750 1.5600 4.7750 0.8300 4.2950 0.8300
                 4.2950 1.3400 3.5950 1.3400 3.5950 1.0900 3.7150 1.0900 3.7150 1.2200 4.1750 1.2200
                 4.1750 0.7100 5.2950 0.7100 5.2950 0.6000 5.5950 0.6000 ;
        POLYGON  4.6550 1.0700 4.5350 1.0700 4.5350 1.5800 4.0950 1.5800 4.0950 1.8700 3.9750 1.8700
                 3.9750 1.5800 3.1950 1.5800 3.1950 1.6100 2.9550 1.6100 2.9550 1.5800 2.4400 1.5800
                 2.4400 1.2900 2.3200 1.2900 2.3200 1.1700 2.5600 1.1700 2.5600 1.4600 3.3550 1.4600
                 3.3550 0.6000 3.6150 0.6000 3.6150 0.7200 3.4750 0.7200 3.4750 1.4600 4.4150 1.4600
                 4.4150 0.9500 4.6550 0.9500 ;
    END
END SDFFRHQX4

MACRO SDFFRHQX2
    CLASS CORE ;
    FOREIGN SDFFRHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2450 1.0900 1.3800 1.5250 ;
        RECT  1.2150 1.0900 1.3800 1.5050 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5650 1.2200 2.8850 1.4100 ;
        RECT  2.5650 1.1800 2.8050 1.4100 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6450 0.9300 7.7650 1.1700 ;
        RECT  7.3200 0.9300 7.7650 1.0500 ;
        RECT  7.3200 0.8850 7.4700 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.9650 1.2550 9.2650 1.4850 ;
        RECT  9.0050 1.2300 9.2650 1.4850 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0050 0.9900 9.5250 1.1100 ;
        RECT  8.1250 0.9700 9.2650 1.0900 ;
        RECT  8.7150 0.9400 8.9750 1.0900 ;
        RECT  8.1250 0.9700 8.2450 1.4400 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5850 1.4650 0.8000 1.7250 ;
        RECT  0.5750 1.3800 0.7700 1.5000 ;
        RECT  0.5850 1.3800 0.7050 2.0300 ;
        RECT  0.5750 0.8000 0.6950 1.5000 ;
        RECT  0.5550 0.6800 0.6750 0.9200 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.1850 -0.1800 9.3050 0.8200 ;
        RECT  7.6450 -0.1800 7.7650 0.6400 ;
        RECT  4.9850 -0.1800 5.2250 0.3900 ;
        RECT  2.7050 0.3800 2.9450 0.5000 ;
        RECT  2.7050 -0.1800 2.8250 0.5000 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  9.0250 1.8450 9.1450 2.7900 ;
        RECT  7.5250 2.2800 7.7650 2.7900 ;
        RECT  5.5850 2.2600 5.8250 2.7900 ;
        RECT  4.7450 2.0100 4.8650 2.7900 ;
        RECT  4.6250 2.0100 4.8650 2.1300 ;
        RECT  3.0050 2.0100 3.1250 2.7900 ;
        RECT  2.8850 2.0100 3.1250 2.1300 ;
        RECT  1.9850 2.0100 2.1050 2.7900 ;
        RECT  1.0050 1.6250 1.1250 2.7900 ;
        RECT  0.1650 1.3800 0.2850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.7650 1.7250 9.6250 1.7250 9.6250 1.8450 9.5050 1.8450 9.5050 1.7250 8.5250 1.7250
                 8.5250 1.2400 8.6450 1.2400 8.6450 1.6050 9.6450 1.6050 9.6450 0.8200 9.6050 0.8200
                 9.6050 0.5800 9.7250 0.5800 9.7250 0.7000 9.7650 0.7000 ;
        POLYGON  8.6650 0.8200 8.0050 0.8200 8.0050 1.5600 8.4050 1.5600 8.4050 2.2100 8.2850 2.2100
                 8.2850 1.6800 8.0050 1.6800 8.0050 1.8000 7.7400 1.8000 7.7400 1.9800 6.8350 1.9800
                 6.8350 1.3000 6.4450 1.3000 6.4450 0.6000 6.7450 0.6000 6.7450 0.7200 6.5650 0.7200
                 6.5650 1.1800 6.9550 1.1800 6.9550 1.8600 7.6200 1.8600 7.6200 1.6800 7.8850 1.6800
                 7.8850 0.7000 8.5450 0.7000 8.5450 0.5600 8.6650 0.5600 ;
        POLYGON  7.4050 1.7400 7.0800 1.7400 7.0800 1.0600 6.6850 1.0600 6.6850 0.9400 6.8650 0.9400
                 6.8650 0.4800 5.9650 0.4800 5.9650 0.8600 6.0850 0.8600 6.0850 1.1000 5.8450 1.1000
                 5.8450 0.6300 4.7450 0.6300 4.7450 0.4800 4.2650 0.4800 4.2650 0.9900 4.4450 0.9900
                 4.4450 1.1100 4.1450 1.1100 4.1450 0.3600 4.8650 0.3600 4.8650 0.5100 5.8450 0.5100
                 5.8450 0.3600 6.9850 0.3600 6.9850 0.5900 7.2000 0.5900 7.2000 1.6200 7.4050 1.6200 ;
        POLYGON  7.4050 2.2200 5.9450 2.2200 5.9450 2.1400 5.2500 2.1400 5.2500 2.0100 4.9850 2.0100
                 4.9850 1.8900 4.2900 1.8900 4.2900 2.2300 3.3250 2.2300 3.3250 1.8900 1.4250 1.8900
                 1.4250 1.6450 1.5000 1.6450 1.5000 0.9200 1.4550 0.9200 1.4550 0.6800 1.5750 0.6800
                 1.5750 0.8000 1.6200 0.8000 1.6200 1.7700 3.3250 1.7700 3.3250 0.8600 3.4450 0.8600
                 3.4450 2.1100 3.9050 2.1100 3.9050 1.1500 4.0250 1.1500 4.0250 2.1100 4.1700 2.1100
                 4.1700 1.7700 5.1050 1.7700 5.1050 1.8900 5.3700 1.8900 5.3700 2.0200 6.0650 2.0200
                 6.0650 2.1000 7.4050 2.1000 ;
        POLYGON  6.5350 1.9400 6.4150 1.9400 6.4150 1.5400 6.2050 1.5400 6.2050 1.3400 4.9250 1.3400
                 4.9250 1.1100 4.8050 1.1100 4.8050 0.9900 5.0450 0.9900 5.0450 1.2200 6.2050 1.2200
                 6.2050 0.7200 6.0850 0.7200 6.0850 0.6000 6.3250 0.6000 6.3250 1.4200 6.5350 1.4200 ;
        POLYGON  6.1150 1.9000 5.9950 1.9000 5.9950 1.7800 5.7300 1.7800 5.7300 1.7700 5.2250 1.7700
                 5.2250 1.6500 5.1050 1.6500 5.1050 1.5300 5.3450 1.5300 5.3450 1.6500 5.8500 1.6500
                 5.8500 1.6600 6.1150 1.6600 ;
        POLYGON  5.7250 1.1000 5.6050 1.1000 5.6050 0.8700 4.6850 0.8700 4.6850 1.6500 4.1450 1.6500
                 4.1450 1.5300 4.5650 1.5300 4.5650 0.8700 4.3850 0.8700 4.3850 0.6000 4.6250 0.6000
                 4.6250 0.7500 5.7250 0.7500 ;
        POLYGON  3.7850 1.9900 3.6650 1.9900 3.6650 0.7400 2.2050 0.7400 2.2050 1.1200 2.0850 1.1200
                 2.0850 0.6200 3.6650 0.6200 3.6650 0.5400 3.7850 0.5400 ;
        POLYGON  3.0850 1.1000 2.9650 1.1000 2.9650 1.0600 2.4450 1.0600 2.4450 1.5300 2.6450 1.5300
                 2.6450 1.6500 2.3250 1.6500 2.3250 1.3600 1.8450 1.3600 1.8450 0.5600 1.3350 0.5600
                 1.3350 0.9700 0.9350 0.9700 0.9350 1.2600 0.8150 1.2600 0.8150 0.8500 1.2150 0.8500
                 1.2150 0.4400 1.9650 0.4400 1.9650 1.2400 2.3250 1.2400 2.3250 0.9400 2.9650 0.9400
                 2.9650 0.8600 3.0850 0.8600 ;
    END
END SDFFRHQX2

MACRO SDFFRHQX1
    CLASS CORE ;
    FOREIGN SDFFRHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1650 0.9150 1.4350 ;
        RECT  0.6500 1.1500 0.8000 1.4350 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3050 1.2300 2.5950 1.3900 ;
        RECT  2.1450 1.1900 2.4250 1.3200 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3050 0.9300 7.4250 1.1700 ;
        RECT  7.0300 0.9300 7.4250 1.0500 ;
        RECT  7.0300 0.8850 7.1800 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4250 1.2100 8.8850 1.3550 ;
        RECT  8.4250 1.2100 8.6850 1.3900 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0450 0.9700 9.1650 1.2100 ;
        RECT  7.7850 0.9700 9.1650 1.0900 ;
        RECT  8.7150 0.9400 8.9750 1.0900 ;
        RECT  7.7850 0.9700 7.9050 1.4400 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 2.0100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.8450 -0.1800 8.9650 0.8200 ;
        RECT  7.3050 -0.1800 7.4250 0.6400 ;
        RECT  4.6250 -0.1800 4.8650 0.3900 ;
        RECT  2.2850 0.3900 2.5250 0.5100 ;
        RECT  2.2850 -0.1800 2.4050 0.5100 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.6850 1.7500 8.8050 2.7900 ;
        RECT  7.2450 2.2200 7.3650 2.7900 ;
        RECT  5.1850 2.2800 5.4250 2.7900 ;
        RECT  4.2250 2.0100 4.3450 2.7900 ;
        RECT  4.1050 2.0100 4.3450 2.1300 ;
        RECT  2.5650 1.7500 2.6850 2.7900 ;
        RECT  2.4450 1.7500 2.6850 1.9300 ;
        RECT  1.3650 2.0100 1.6050 2.1300 ;
        RECT  1.3650 2.0100 1.4850 2.7900 ;
        RECT  0.5550 1.5550 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.4050 1.6800 9.3250 1.6800 9.3250 1.8000 9.2050 1.8000 9.2050 1.6300 8.1850 1.6300
                 8.1850 1.2400 8.3050 1.2400 8.3050 1.5100 9.2850 1.5100 9.2850 0.8500 9.2650 0.8500
                 9.2650 0.5800 9.3850 0.5800 9.3850 0.7300 9.4050 0.7300 ;
        POLYGON  8.3250 0.8500 7.6650 0.8500 7.6650 1.5600 8.0650 1.5600 8.0650 2.2100 7.9450 2.2100
                 7.9450 1.6800 7.6650 1.6800 7.6650 1.9800 6.4750 1.9800 6.4750 1.3000 6.0150 1.3000
                 6.0150 0.7200 5.9650 0.7200 5.9650 0.6000 6.2050 0.6000 6.2050 0.7200 6.1350 0.7200
                 6.1350 1.1800 6.5950 1.1800 6.5950 1.8600 7.5450 1.8600 7.5450 0.7300 8.2050 0.7300
                 8.2050 0.5900 8.3250 0.5900 ;
        POLYGON  7.1050 2.2200 5.5450 2.2200 5.5450 2.1600 4.4650 2.1600 4.4650 1.8900 3.5050 1.8900
                 3.5050 2.2300 2.9050 2.2300 2.9050 1.6300 2.3250 1.6300 2.3250 1.8900 0.9750 1.8900
                 0.9750 1.5550 1.0350 1.5550 1.0350 0.6800 1.1550 0.6800 1.1550 1.7700 2.2050 1.7700
                 2.2050 1.5100 2.9050 1.5100 2.9050 0.8700 3.0250 0.8700 3.0250 2.1100 3.3850 2.1100
                 3.3850 1.2700 3.4850 1.2700 3.4850 1.1500 3.6050 1.1500 3.6050 1.3900 3.5050 1.3900
                 3.5050 1.7700 4.5850 1.7700 4.5850 2.0400 5.6650 2.0400 5.6650 2.1000 7.1050 2.1000 ;
        POLYGON  7.0450 1.7400 6.7900 1.7400 6.7900 1.0600 6.2550 1.0600 6.2550 0.9400 6.3750 0.9400
                 6.3750 0.4800 5.4250 0.4800 5.4250 0.8600 5.5850 0.8600 5.5850 1.1000 5.3050 1.1000
                 5.3050 0.6300 4.3850 0.6300 4.3850 0.4800 3.9050 0.4800 3.9050 0.9200 4.0250 0.9200
                 4.0250 1.0400 3.7850 1.0400 3.7850 0.3600 4.5050 0.3600 4.5050 0.5100 5.3050 0.5100
                 5.3050 0.3600 6.4950 0.3600 6.4950 0.9400 6.7900 0.9400 6.7900 0.5900 6.9100 0.5900
                 6.9100 1.6200 7.0450 1.6200 ;
        POLYGON  6.1750 1.9400 6.0550 1.9400 6.0550 1.5400 5.8250 1.5400 5.8250 1.5600 4.5050 1.5600
                 4.5050 1.1100 4.3850 1.1100 4.3850 0.9900 4.6250 0.9900 4.6250 1.4400 5.7050 1.4400
                 5.7050 0.7200 5.5450 0.7200 5.5450 0.6000 5.8250 0.6000 5.8250 1.4200 6.1750 1.4200 ;
        POLYGON  5.7550 1.9200 4.7050 1.9200 4.7050 1.6800 4.9450 1.6800 4.9450 1.8000 5.6350 1.8000
                 5.6350 1.6800 5.7550 1.6800 ;
        POLYGON  5.1450 1.3200 5.0250 1.3200 5.0250 0.8700 4.2650 0.8700 4.2650 1.6500 3.6250 1.6500
                 3.6250 1.5300 4.1450 1.5300 4.1450 0.7200 4.0250 0.7200 4.0250 0.6000 4.2650 0.6000
                 4.2650 0.7500 5.1450 0.7500 ;
        POLYGON  3.2650 1.9900 3.1450 1.9900 3.1450 0.7500 1.7850 0.7500 1.7850 1.1200 1.6650 1.1200
                 1.6650 0.6300 3.1450 0.6300 3.1450 0.5400 3.2650 0.5400 ;
        POLYGON  2.6650 1.1100 2.5450 1.1100 2.5450 1.0700 2.0250 1.0700 2.0250 1.5300 2.0850 1.5300
                 2.0850 1.6500 1.8450 1.6500 1.8450 1.5300 1.9050 1.5300 1.9050 1.3600 1.4250 1.3600
                 1.4250 0.5600 0.9150 0.5600 0.9150 1.0300 0.5150 1.0300 0.5150 1.2600 0.3950 1.2600
                 0.3950 0.9100 0.7950 0.9100 0.7950 0.4400 1.5450 0.4400 1.5450 1.2400 1.9050 1.2400
                 1.9050 0.9500 2.5450 0.9500 2.5450 0.8700 2.6650 0.8700 ;
    END
END SDFFRHQX1

MACRO SDFFQXL
    CLASS CORE ;
    FOREIGN SDFFQXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.3200 0.8950 1.6250 ;
        RECT  0.6500 1.4100 0.8000 1.7250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2350 1.2300 5.8650 1.3500 ;
        RECT  5.2350 1.2300 5.4950 1.3800 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6850 1.2450 7.1850 1.3900 ;
        RECT  6.6850 1.2100 6.9450 1.3900 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4450 0.9500 7.4450 1.0700 ;
        RECT  6.9750 0.9400 7.2350 1.0900 ;
        RECT  6.5850 0.9400 7.2350 1.0700 ;
        RECT  6.5850 0.9300 6.8250 1.0700 ;
        RECT  6.4450 0.9500 6.5650 1.3900 ;
        RECT  6.2250 1.4700 6.4650 1.5900 ;
        RECT  6.3450 1.2700 6.4650 1.5900 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1950 1.3200 0.3150 1.9650 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4400 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  7.1450 -0.1800 7.2650 0.7900 ;
        RECT  5.8650 -0.1800 5.9850 0.7900 ;
        RECT  3.6950 -0.1800 3.9350 0.3400 ;
        RECT  2.0150 -0.1800 2.2550 0.3400 ;
        RECT  0.5550 -0.1800 0.6750 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  7.0850 1.9500 7.3250 2.0700 ;
        RECT  7.0850 1.9500 7.2050 2.7900 ;
        RECT  5.7250 1.9500 5.9650 2.0700 ;
        RECT  5.7250 1.9500 5.8450 2.7900 ;
        RECT  3.6950 2.0800 3.9350 2.2000 ;
        RECT  3.6950 2.0800 3.8150 2.7900 ;
        RECT  2.0950 2.0800 2.3350 2.2000 ;
        RECT  2.0950 2.0800 2.2150 2.7900 ;
        RECT  0.6150 1.8450 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.6850 2.0100 7.5650 2.0100 7.5650 1.6300 6.5850 1.6300 6.5850 1.5100 7.5650 1.5100
                 7.5650 0.5500 7.6850 0.5500 ;
        POLYGON  6.6250 0.8100 6.3250 0.8100 6.3250 1.1500 6.1050 1.1500 6.1050 1.7100 6.4650 1.7100
                 6.4650 1.7700 6.5450 1.7700 6.5450 2.0100 6.4250 2.0100 6.4250 1.8900 6.3450 1.8900
                 6.3450 1.8300 4.9350 1.8300 4.9350 1.5900 4.9950 1.5900 4.9950 0.7400 5.2350 0.7400
                 5.2350 0.8600 5.1150 0.8600 5.1150 1.7100 5.9850 1.7100 5.9850 1.0300 6.2050 1.0300
                 6.2050 0.6900 6.5050 0.6900 6.5050 0.5500 6.6250 0.5500 ;
        POLYGON  5.6250 0.7300 5.3850 0.7300 5.3850 0.6200 4.8750 0.6200 4.8750 1.4600 4.8150 1.4600
                 4.8150 1.9500 5.5450 1.9500 5.5450 2.0700 4.6950 2.0700 4.6950 1.2200 4.7550 1.2200
                 4.7550 0.6200 3.1950 0.6200 3.1950 1.2400 3.0750 1.2400 3.0750 0.5000 4.2550 0.5000
                 4.2550 0.4200 4.4950 0.4200 4.4950 0.5000 5.5050 0.5000 5.5050 0.6100 5.6250 0.6100 ;
        POLYGON  4.6350 0.8600 4.5150 0.8600 4.5150 1.3800 4.5750 1.3800 4.5750 1.7800 4.4550 1.7800
                 4.4550 1.5000 3.7350 1.5000 3.7350 1.3800 3.5750 1.3800 3.5750 1.2600 3.8550 1.2600
                 3.8550 1.3800 4.3950 1.3800 4.3950 0.7400 4.6350 0.7400 ;
        POLYGON  4.4950 2.1600 4.2550 2.1600 4.2550 2.0200 4.0650 2.0200 4.0650 1.9600 3.3900 1.9600
                 3.3900 2.0200 3.1750 2.0200 3.1750 2.1600 2.9350 2.1600 2.9350 2.0200 2.4750 2.0200
                 2.4750 1.9600 1.1550 1.9600 1.1550 1.9650 1.0350 1.9650 1.0350 0.7400 1.2750 0.7400
                 1.2750 0.8600 1.1550 0.8600 1.1550 1.8400 2.4750 1.8400 2.4750 1.0600 2.7150 1.0600
                 2.7150 1.1800 2.5950 1.1800 2.5950 1.9000 3.2700 1.9000 3.2700 1.8400 4.1850 1.8400
                 4.1850 1.9000 4.3750 1.9000 4.3750 2.0400 4.4950 2.0400 ;
        POLYGON  4.0950 1.2600 3.9750 1.2600 3.9750 1.1400 3.4550 1.1400 3.4550 1.7200 3.2150 1.7200
                 3.2150 1.6000 3.3350 1.6000 3.3350 0.8600 3.3150 0.8600 3.3150 0.7400 3.5550 0.7400
                 3.5550 0.8600 3.4550 0.8600 3.4550 1.0200 4.0950 1.0200 ;
        POLYGON  2.9750 1.7800 2.8550 1.7800 2.8550 1.4800 2.8350 1.4800 2.8350 0.9200 2.6750 0.9200
                 2.6750 0.6800 2.3050 0.6800 2.3050 0.5800 1.7750 0.5800 1.7750 0.5200 1.6350 0.5200
                 1.6350 0.4000 1.8950 0.4000 1.8950 0.4600 2.4250 0.4600 2.4250 0.5600 2.7950 0.5600
                 2.7950 0.8000 2.9550 0.8000 2.9550 1.3600 2.9750 1.3600 ;
        POLYGON  2.3550 1.2600 1.7350 1.2600 1.7350 1.6000 1.8550 1.6000 1.8550 1.7200 1.6150 1.7200
                 1.6150 0.9200 1.5350 0.9200 1.5350 0.8000 1.3950 0.8000 1.3950 0.6200 0.9150 0.6200
                 0.9150 1.2000 0.3950 1.2000 0.3950 1.0800 0.7950 1.0800 0.7950 0.5000 1.5150 0.5000
                 1.5150 0.6800 1.6550 0.6800 1.6550 0.8000 1.7350 0.8000 1.7350 1.1400 2.3550 1.1400 ;
    END
END SDFFQXL

MACRO SDFFQX4
    CLASS CORE ;
    FOREIGN SDFFQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9150 0.7200 2.1550 0.8400 ;
        RECT  1.9350 1.2800 2.0550 2.0400 ;
        RECT  1.9150 0.7200 2.0350 1.4000 ;
        RECT  0.9400 1.0250 2.0350 1.1450 ;
        RECT  1.0950 0.7200 1.2150 2.0400 ;
        RECT  0.9400 0.8850 1.2150 1.1450 ;
        RECT  0.9550 0.7200 1.2150 1.1450 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4750 0.9800 0.8000 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        RECT  0.4750 0.9800 0.5950 1.2200 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.1600 7.5250 1.3800 ;
        RECT  7.3850 1.1200 7.5050 1.5100 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4250 1.2200 8.7450 1.4400 ;
        RECT  8.4250 1.2200 8.6850 1.4650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8850 0.9800 9.0650 1.1000 ;
        RECT  8.7150 0.9400 8.9750 1.1000 ;
        RECT  7.6450 1.3900 8.0050 1.5100 ;
        RECT  7.8850 0.9800 8.0050 1.5100 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.7250 -0.1800 8.8450 0.8200 ;
        RECT  7.2650 0.6400 7.5050 0.7600 ;
        RECT  7.3850 -0.1800 7.5050 0.7600 ;
        RECT  5.1750 -0.1800 5.2950 0.3800 ;
        RECT  3.4750 -0.1800 3.5950 0.3800 ;
        RECT  2.3950 -0.1800 2.6350 0.3600 ;
        RECT  1.4350 -0.1800 1.6750 0.3600 ;
        RECT  0.4750 -0.1800 0.5950 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.5650 1.9300 8.8050 2.0500 ;
        RECT  8.5650 1.9300 8.6850 2.7900 ;
        RECT  7.2250 1.8700 7.3450 2.7900 ;
        RECT  4.9350 2.2000 5.1750 2.7900 ;
        RECT  3.2550 1.6600 3.3750 2.7900 ;
        RECT  2.3550 1.3900 2.4750 2.7900 ;
        RECT  1.5150 1.3900 1.6350 2.7900 ;
        RECT  0.6750 1.3900 0.7950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.3050 1.8250 9.1650 1.8250 9.1650 1.9900 9.0450 1.9900 9.0450 1.7050 8.1250 1.7050
                 8.1250 1.4300 8.2450 1.4300 8.2450 1.5850 9.1850 1.5850 9.1850 0.8200 9.1450 0.8200
                 9.1450 0.5800 9.2650 0.5800 9.2650 0.7000 9.3050 0.7000 ;
        POLYGON  8.2050 0.8200 7.7650 0.8200 7.7650 1.0000 7.1450 1.0000 7.1450 1.6300 7.9850 1.6300
                 7.9850 1.9900 7.8650 1.9900 7.8650 1.7500 6.3750 1.7500 6.3750 1.9000 6.2550 1.9000
                 6.2550 1.6300 7.0250 1.6300 7.0250 0.5200 6.5150 0.5200 6.5150 0.8400 6.2750 0.8400
                 6.2750 0.7200 6.3950 0.7200 6.3950 0.4000 7.1450 0.4000 7.1450 0.8800 7.6450 0.8800
                 7.6450 0.7000 8.0850 0.7000 8.0850 0.5800 8.2050 0.5800 ;
        POLYGON  6.9850 2.0500 6.8650 2.0500 6.8650 2.1400 6.0150 2.1400 6.0150 2.0800 4.2150 2.0800
                 4.2150 1.4400 4.0350 1.4400 4.0350 1.5600 3.9150 1.5600 3.9150 1.3200 4.2150 1.3200
                 4.2150 1.1200 4.4550 1.1200 4.4550 1.0000 4.5750 1.0000 4.5750 1.2400 4.3350 1.2400
                 4.3350 1.9600 6.0150 1.9600 6.0150 1.3200 6.6350 1.3200 6.6350 0.6400 6.9050 0.6400
                 6.9050 0.7600 6.7550 0.7600 6.7550 1.4400 6.1350 1.4400 6.1350 2.0200 6.7450 2.0200
                 6.7450 1.9300 6.9850 1.9300 ;
        POLYGON  6.2750 1.1600 6.0350 1.1600 6.0350 0.5400 5.6750 0.5400 5.6750 0.6200 5.6550 0.6200
                 5.6550 1.5600 5.5350 1.5600 5.5350 0.6200 4.9350 0.6200 4.9350 0.5400 3.8550 0.5400
                 3.8550 0.6200 3.2350 0.6200 3.2350 0.6000 0.8350 0.6000 0.8350 0.6600 0.2550 0.6600
                 0.2550 1.3900 0.3150 1.3900 0.3150 1.6300 0.1950 1.6300 0.1950 1.5100 0.1350 1.5100
                 0.1350 0.5400 0.7150 0.5400 0.7150 0.4800 3.3550 0.4800 3.3550 0.5000 3.7350 0.5000
                 3.7350 0.4200 3.9350 0.4200 3.9350 0.4000 4.1750 0.4000 4.1750 0.4200 5.0550 0.4200
                 5.0550 0.5000 5.5550 0.5000 5.5550 0.4200 6.1550 0.4200 6.1550 1.0400 6.2750 1.0400 ;
        POLYGON  5.9150 1.2000 5.8950 1.2000 5.8950 1.8400 5.6550 1.8400 5.6550 1.8000 5.2950 1.8000
                 5.2950 1.5000 4.9350 1.5000 4.9350 1.3800 5.4150 1.3800 5.4150 1.6800 5.7750 1.6800
                 5.7750 1.0800 5.7950 1.0800 5.7950 0.6600 5.9150 0.6600 ;
        POLYGON  5.3150 1.2200 5.1950 1.2200 5.1950 1.1000 4.8150 1.1000 4.8150 1.8400 4.4550 1.8400
                 4.4550 1.7200 4.6950 1.7200 4.6950 0.6600 4.8150 0.6600 4.8150 0.9800 5.3150 0.9800 ;
        POLYGON  4.4550 0.8400 4.0950 0.8400 4.0950 1.2000 3.7950 1.2000 3.7950 1.6800 3.9750 1.6800
                 3.9750 1.7200 4.0950 1.7200 4.0950 1.8400 3.8550 1.8400 3.8550 1.8000 3.6750 1.8000
                 3.6750 1.4600 3.0750 1.4600 3.0750 1.2000 3.1950 1.2000 3.1950 1.3400 3.6750 1.3400
                 3.6750 1.0800 3.9750 1.0800 3.9750 0.7200 4.4550 0.7200 ;
        POLYGON  3.5550 1.2200 3.4350 1.2200 3.4350 1.0800 2.9550 1.0800 2.9550 2.0400 2.8350 2.0400
                 2.8350 1.0800 2.3950 1.0800 2.3950 1.1600 2.1550 1.1600 2.1550 0.9600 2.8350 0.9600
                 2.8350 0.7200 3.1150 0.7200 3.1150 0.8400 2.9550 0.8400 2.9550 0.9600 3.5550 0.9600 ;
    END
END SDFFQX4

MACRO SDFFQX2
    CLASS CORE ;
    FOREIGN SDFFQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.0900 1.3800 1.5900 ;
        RECT  1.2300 1.0900 1.3800 1.5600 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8700 1.1900 6.1800 1.4300 ;
        RECT  5.8700 1.1750 6.0200 1.4350 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5550 1.2100 7.8150 1.4100 ;
        RECT  7.3400 1.2100 7.8150 1.3800 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7400 0.9700 7.9000 1.0900 ;
        RECT  7.0800 0.9400 7.5250 1.0900 ;
        RECT  7.0800 0.9100 7.2000 1.1500 ;
        RECT  6.5400 1.2300 6.8600 1.3500 ;
        RECT  6.7400 0.9700 6.8600 1.3500 ;
        RECT  6.5400 1.2300 6.6600 1.4700 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6000 0.6800 0.7200 2.0400 ;
        RECT  0.3600 0.8850 0.7200 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.5600 -0.1800 7.6800 0.7900 ;
        RECT  6.2600 -0.1800 6.3800 0.7900 ;
        RECT  4.1300 -0.1800 4.3700 0.3700 ;
        RECT  2.2500 0.6300 2.4900 0.7500 ;
        RECT  2.2500 -0.1800 2.3700 0.7500 ;
        RECT  1.0200 -0.1800 1.1400 0.7300 ;
        RECT  0.1800 -0.1800 0.3000 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.4400 1.9100 7.5600 2.7900 ;
        RECT  6.1600 1.9100 6.2800 2.7900 ;
        RECT  4.1100 2.2300 4.2300 2.7900 ;
        RECT  2.2700 2.0100 2.5100 2.1300 ;
        RECT  2.2700 2.0100 2.3900 2.7900 ;
        RECT  1.0200 1.6800 1.1400 2.7900 ;
        RECT  0.1800 1.3900 0.3000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.1400 1.7700 7.9800 1.7700 7.9800 2.0300 7.8600 2.0300 7.8600 1.6500 7.1000 1.6500
                 7.1000 1.4300 6.9800 1.4300 6.9800 1.3100 7.2200 1.3100 7.2200 1.5300 8.0200 1.5300
                 8.0200 0.7900 7.9800 0.7900 7.9800 0.5500 8.1000 0.5500 8.1000 0.6700 8.1400 0.6700 ;
        POLYGON  7.0400 0.7900 6.6200 0.7900 6.6200 1.1100 6.4200 1.1100 6.4200 1.5900 6.9200 1.5900
                 6.9200 2.0300 6.8000 2.0300 6.8000 1.7100 5.6100 1.7100 5.6100 1.8100 5.2900 1.8100
                 5.2900 1.6900 5.4900 1.6900 5.4900 0.9100 5.4300 0.9100 5.4300 0.6700 5.5500 0.6700
                 5.5500 0.7900 5.6100 0.7900 5.6100 1.5900 6.3000 1.5900 6.3000 0.9900 6.5000 0.9900
                 6.5000 0.6700 6.9200 0.6700 6.9200 0.5500 7.0400 0.5500 ;
        POLYGON  5.9600 0.7900 5.8400 0.7900 5.8400 0.5500 5.3100 0.5500 5.3100 1.0900 5.1700 1.0900
                 5.1700 1.3700 5.3700 1.3700 5.3700 1.4900 5.1700 1.4900 5.1700 1.9300 5.9200 1.9300
                 5.9200 2.0500 5.0500 2.0500 5.0500 0.9700 5.1900 0.9700 5.1900 0.5500 4.6100 0.5500
                 4.6100 0.6100 3.5300 0.6100 3.5300 1.2300 3.4100 1.2300 3.4100 0.4900 4.4900 0.4900
                 4.4900 0.4300 4.6900 0.4300 4.6900 0.4100 4.9300 0.4100 4.9300 0.4300 5.9600 0.4300 ;
        POLYGON  5.0700 0.8500 4.9300 0.8500 4.9300 1.8700 4.8100 1.8700 4.8100 1.4900 3.8900 1.4900
                 3.8900 1.3700 4.8100 1.3700 4.8100 0.7300 5.0700 0.7300 ;
        POLYGON  4.8500 2.2500 4.3500 2.2500 4.3500 2.1100 3.5300 2.1100 3.5300 2.2500 3.2900 2.2500
                 3.2900 2.1100 2.8300 2.1100 2.8300 1.8900 1.5600 1.8900 1.5600 1.9500 1.4400 1.9500
                 1.4400 1.7100 1.5000 1.7100 1.5000 0.6800 1.6200 0.6800 1.6200 1.7700 2.8300 1.7700
                 2.8300 1.2300 2.8100 1.2300 2.8100 1.1100 3.0500 1.1100 3.0500 1.2300 2.9500 1.2300
                 2.9500 1.9900 4.4700 1.9900 4.4700 2.1300 4.8500 2.1300 ;
        POLYGON  4.4900 1.2500 3.7700 1.2500 3.7700 1.7500 3.7500 1.7500 3.7500 1.8700 3.6300 1.8700
                 3.6300 1.6300 3.6500 1.6300 3.6500 0.7300 3.8900 0.7300 3.8900 0.8500 3.7700 0.8500
                 3.7700 1.1300 4.4900 1.1300 ;
        POLYGON  3.3300 1.8700 3.2100 1.8700 3.2100 1.4700 3.1700 1.4700 3.1700 0.9100 2.8200 0.9100
                 2.8200 0.9900 2.2900 0.9900 2.2900 1.2300 2.1700 1.2300 2.1700 0.8700 2.7000 0.8700
                 2.7000 0.7900 3.1300 0.7900 3.1300 0.6700 3.2500 0.6700 3.2500 0.7900 3.2900 0.7900
                 3.2900 1.3500 3.3300 1.3500 ;
        POLYGON  2.7100 1.4700 2.0300 1.4700 2.0300 1.6500 1.7900 1.6500 1.7900 1.5300 1.9100 1.5300
                 1.9100 0.9100 1.8900 0.9100 1.8900 0.6700 1.7900 0.6700 1.7900 0.5600 1.3800 0.5600
                 1.3800 0.9700 1.0000 0.9700 1.0000 1.2400 0.8800 1.2400 0.8800 0.8500 1.2600 0.8500
                 1.2600 0.4400 1.9100 0.4400 1.9100 0.5500 2.0100 0.5500 2.0100 0.7900 2.0300 0.7900
                 2.0300 1.3500 2.7100 1.3500 ;
    END
END SDFFQX2

MACRO SDFFQX1
    CLASS CORE ;
    FOREIGN SDFFQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.2200 0.8950 1.4600 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.3400 0.8000 1.7250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6050 1.2100 5.7250 1.4500 ;
        RECT  5.2350 1.2300 5.7250 1.3800 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6850 1.2100 7.0450 1.4100 ;
        RECT  6.6850 1.2100 6.9450 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.2050 0.8900 7.3450 1.0100 ;
        RECT  6.9750 0.8900 7.2350 1.0900 ;
        RECT  6.5050 0.7700 6.6250 1.0100 ;
        RECT  6.2050 0.8900 6.3250 1.4300 ;
        RECT  6.0850 1.3100 6.2050 1.5500 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 2.2100 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  7.0050 1.9700 7.1250 2.7900 ;
        RECT  5.7250 1.9700 5.8450 2.7900 ;
        RECT  3.6750 2.2000 3.7950 2.7900 ;
        RECT  2.0150 2.1400 2.2550 2.2600 ;
        RECT  2.0150 2.1400 2.1350 2.7900 ;
        RECT  0.5550 1.8450 0.6750 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  7.0050 -0.1800 7.1250 0.6500 ;
        RECT  5.7250 -0.1800 5.8450 0.6500 ;
        RECT  3.6150 -0.1800 3.8550 0.3400 ;
        RECT  1.8750 -0.1800 2.1150 0.3200 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  7.5850 1.7950 7.5450 1.7950 7.5450 2.0900 7.4250 2.0900 7.4250 1.6750 6.4450 1.6750
                 6.4450 1.1300 6.5650 1.1300 6.5650 1.5550 7.4650 1.5550 7.4650 0.7700 7.4250 0.7700
                 7.4250 0.4100 7.5450 0.4100 7.5450 0.6500 7.5850 0.6500 ;
        POLYGON  6.4850 0.6500 6.0850 0.6500 6.0850 1.1900 5.9650 1.1900 5.9650 1.6700 6.3250 1.6700
                 6.3250 1.7950 6.4850 1.7950 6.4850 2.0900 6.3650 2.0900 6.3650 1.9150 6.2050 1.9150
                 6.2050 1.7900 4.8550 1.7900 4.8550 1.6700 4.9150 1.6700 4.9150 0.6800 5.0350 0.6800
                 5.0350 1.6700 5.8450 1.6700 5.8450 1.0700 5.9650 1.0700 5.9650 0.5300 6.3650 0.5300
                 6.3650 0.4100 6.4850 0.4100 ;
        POLYGON  5.4850 2.0300 4.6150 2.0300 4.6150 1.2800 4.6750 1.2800 4.6750 0.5600 4.1750 0.5600
                 4.1750 0.5800 3.1150 0.5800 3.1150 1.2400 2.9950 1.2400 2.9950 0.4600 4.0550 0.4600
                 4.0550 0.4400 4.1550 0.4400 4.1550 0.4000 4.3950 0.4000 4.3950 0.4400 5.3050 0.4400
                 5.3050 0.4100 5.4250 0.4100 5.4250 0.6500 5.3050 0.6500 5.3050 0.5600 4.7950 0.5600
                 4.7950 1.5200 4.7350 1.5200 4.7350 1.9100 5.4850 1.9100 ;
        POLYGON  4.5550 0.8600 4.4950 0.8600 4.4950 1.8400 4.3750 1.8400 4.3750 1.4400 3.4950 1.4400
                 3.4950 1.3200 4.3750 1.3200 4.3750 0.8600 4.3150 0.8600 4.3150 0.7400 4.5550 0.7400 ;
        POLYGON  4.4150 2.2200 3.9850 2.2200 3.9850 2.0800 3.1650 2.0800 3.1650 2.2200 2.9250 2.2200
                 2.9250 2.0800 2.3950 2.0800 2.3950 2.0200 1.0350 2.0200 1.0350 0.6800 1.1550 0.6800
                 1.1550 1.9000 2.3950 1.9000 2.3950 1.0600 2.6350 1.0600 2.6350 1.1800 2.5150 1.1800
                 2.5150 1.9600 4.1050 1.9600 4.1050 2.1000 4.4150 2.1000 ;
        POLYGON  4.0750 1.2000 3.3550 1.2000 3.3550 1.7200 3.3150 1.7200 3.3150 1.8400 3.1950 1.8400
                 3.1950 1.6000 3.2350 1.6000 3.2350 0.7400 3.4750 0.7400 3.4750 0.8600 3.3550 0.8600
                 3.3550 1.0800 4.0750 1.0800 ;
        POLYGON  2.8950 1.8400 2.7750 1.8400 2.7750 1.4800 2.7550 1.4800 2.7550 0.9200 2.7150 0.9200
                 2.7150 0.6800 1.6650 0.6800 1.6650 0.5600 1.5150 0.5600 1.5150 0.4000 1.7550 0.4000
                 1.7550 0.4400 1.7850 0.4400 1.7850 0.5600 2.8350 0.5600 2.8350 0.8000 2.8750 0.8000
                 2.8750 1.3600 2.8950 1.3600 ;
        POLYGON  2.2750 1.2600 1.6550 1.2600 1.6550 1.6600 1.7750 1.6600 1.7750 1.7800 1.5350 1.7800
                 1.5350 0.9200 1.4250 0.9200 1.4250 0.8000 1.2750 0.8000 1.2750 0.5600 0.9150 0.5600
                 0.9150 1.1000 0.5350 1.1000 0.5350 1.2400 0.4150 1.2400 0.4150 0.9800 0.7950 0.9800
                 0.7950 0.4400 1.3950 0.4400 1.3950 0.6800 1.5450 0.6800 1.5450 0.8000 1.6550 0.8000
                 1.6550 1.1400 2.2750 1.1400 ;
    END
END SDFFQX1

MACRO SDFFNSRXL
    CLASS CORE ;
    FOREIGN SDFFNSRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.0500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.2300 2.3050 1.5000 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8550 2.1100 7.6350 2.2300 ;
        RECT  6.8550 1.7800 6.9750 2.2300 ;
        RECT  4.4150 1.8800 6.9750 1.9000 ;
        RECT  5.6550 1.7800 6.9750 1.9000 ;
        RECT  5.1750 1.8800 5.7750 2.0000 ;
        RECT  3.3550 1.7800 5.2950 1.8900 ;
        RECT  3.2450 1.7700 4.5350 1.8250 ;
        RECT  3.2450 1.7050 3.4750 1.8250 ;
        RECT  3.2450 1.4650 3.4100 1.8250 ;
        RECT  3.2450 0.9400 3.3650 1.8250 ;
        END
    END SN
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.2150 1.2800 10.4550 1.4000 ;
        RECT  10.1650 1.5200 10.4250 1.6700 ;
        RECT  10.2150 1.2800 10.3350 1.6700 ;
        END
    END CKN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7450 1.5200 11.0050 1.6700 ;
        RECT  10.7550 1.2900 10.9950 1.6700 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 1.4700 12.4550 1.6700 ;
        RECT  11.9650 1.4700 12.4550 1.6350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 0.9400 12.4550 1.0900 ;
        RECT  12.2650 0.9400 12.3850 1.2400 ;
        RECT  11.3650 1.0000 12.3850 1.1200 ;
        RECT  11.4550 0.9600 11.5750 1.2000 ;
        RECT  11.3650 1.0000 11.4850 1.7700 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 0.6800 0.2650 1.5800 ;
        RECT  0.0700 0.8850 0.2650 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4350 1.5100 1.5550 1.7500 ;
        RECT  1.3750 0.6300 1.4950 0.8700 ;
        RECT  1.2300 1.4650 1.4550 1.7250 ;
        RECT  1.3350 0.7500 1.4550 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.0500 0.1800 ;
        RECT  11.9550 -0.1800 12.0750 0.8800 ;
        RECT  10.6750 -0.1800 10.7950 0.8800 ;
        RECT  9.6850 -0.1800 9.9250 0.3400 ;
        RECT  7.8150 -0.1800 7.9350 0.8600 ;
        RECT  3.0850 -0.1800 3.3250 0.3200 ;
        RECT  1.7950 -0.1800 1.9150 0.8700 ;
        RECT  0.5650 -0.1800 0.6850 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.0500 2.7900 ;
        RECT  12.2450 2.0300 12.3650 2.7900 ;
        RECT  10.6750 1.9700 10.7950 2.7900 ;
        RECT  9.8650 2.1200 9.9850 2.7900 ;
        RECT  7.7550 2.2900 7.9950 2.7900 ;
        RECT  6.1350 2.2600 6.3750 2.7900 ;
        RECT  4.4550 2.2600 4.6950 2.7900 ;
        RECT  3.1350 2.2500 3.3750 2.7900 ;
        RECT  1.8550 1.6300 1.9750 2.7900 ;
        RECT  0.5650 1.4600 0.6850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.8450 2.0900 12.7250 2.0900 12.7250 1.9700 12.5750 1.9700 12.5750 1.9100
                 11.7050 1.9100 11.7050 1.5100 11.8250 1.5100 11.8250 1.7900 12.5750 1.7900
                 12.5750 0.8200 12.3450 0.8200 12.3450 0.7000 12.6950 0.7000 12.6950 1.8500
                 12.8450 1.8500 ;
        POLYGON  11.6250 2.1500 11.3850 2.1500 11.3850 2.0300 11.1250 2.0300 11.1250 1.1200
                 10.4350 1.1200 10.4350 0.5800 8.9950 0.5800 8.9950 0.7400 9.0850 0.7400 9.0850 1.3000
                 9.1750 1.3000 9.1750 1.8600 9.2950 1.8600 9.2950 1.9800 9.0550 1.9800 9.0550 1.4200
                 8.9650 1.4200 8.9650 0.8600 8.8750 0.8600 8.8750 0.4600 10.5550 0.4600 10.5550 1.0000
                 11.1250 1.0000 11.1250 0.7600 11.2150 0.7600 11.2150 0.7000 11.4950 0.7000
                 11.4950 0.8200 11.3350 0.8200 11.3350 0.8800 11.2450 0.8800 11.2450 1.9100
                 11.5050 1.9100 11.5050 2.0300 11.6250 2.0300 ;
        POLYGON  10.4350 2.0300 10.1950 2.0300 10.1950 2.0000 9.9250 2.0000 9.9250 1.1600 9.5350 1.1600
                 9.5350 1.0400 10.0750 1.0400 10.0750 0.7000 10.3150 0.7000 10.3150 0.8200
                 10.1950 0.8200 10.1950 1.1600 10.0450 1.1600 10.0450 1.8800 10.4350 1.8800 ;
        POLYGON  9.6250 2.2200 8.2150 2.2200 8.2150 2.1400 7.7550 2.1400 7.7550 1.9900 7.0950 1.9900
                 7.0950 1.6500 6.6950 1.6500 6.6950 1.3600 6.4050 1.3600 6.4050 1.2400 6.8150 1.2400
                 6.8150 1.5300 7.2150 1.5300 7.2150 1.8700 7.8750 1.8700 7.8750 2.0200 8.3350 2.0200
                 8.3350 2.1000 8.8150 2.1000 8.8150 1.6600 8.5150 1.6600 8.5150 1.5400 8.6350 1.5400
                 8.6350 1.1200 8.6050 1.1200 8.6050 1.0000 8.8450 1.0000 8.8450 1.1200 8.7550 1.1200
                 8.7550 1.5400 8.9350 1.5400 8.9350 2.1000 9.5050 2.1000 9.5050 1.6000 9.2950 1.6000
                 9.2950 0.8200 9.2050 0.8200 9.2050 0.7000 9.4450 0.7000 9.4450 0.8200 9.4150 0.8200
                 9.4150 1.4800 9.6250 1.4800 ;
        POLYGON  8.6950 1.9800 8.4550 1.9800 8.4550 1.9000 8.2750 1.9000 8.2750 1.1600 7.1750 1.1600
                 7.1750 1.0400 8.3650 1.0400 8.3650 0.7400 8.4550 0.7400 8.4550 0.6200 8.5750 0.6200
                 8.5750 0.8600 8.4850 0.8600 8.4850 1.1600 8.3950 1.1600 8.3950 1.7800 8.5750 1.7800
                 8.5750 1.8600 8.6950 1.8600 ;
        POLYGON  8.1550 1.4100 7.4550 1.4100 7.4550 1.6300 7.5750 1.6300 7.5750 1.7500 7.3350 1.7500
                 7.3350 1.4100 6.9350 1.4100 6.9350 1.0400 6.2850 1.0400 6.2850 1.6600 5.8850 1.6600
                 5.8850 1.5400 6.1650 1.5400 6.1650 0.6200 6.2850 0.6200 6.2850 0.9200 6.9350 0.9200
                 6.9350 0.8000 6.9750 0.8000 6.9750 0.6200 7.0950 0.6200 7.0950 0.9200 7.0550 0.9200
                 7.0550 1.2900 8.1550 1.2900 ;
        POLYGON  7.5150 0.8600 7.3950 0.8600 7.3950 0.6200 7.2150 0.6200 7.2150 0.5000 6.7350 0.5000
                 6.7350 0.8000 6.4950 0.8000 6.4950 0.6800 6.6150 0.6800 6.6150 0.3800 7.3350 0.3800
                 7.3350 0.5000 7.5150 0.5000 ;
        POLYGON  6.7350 2.1900 6.4950 2.1900 6.4950 2.1400 6.0150 2.1400 6.0150 2.2400 4.9250 2.2400
                 4.9250 2.1400 4.2950 2.1400 4.2950 2.2500 4.1750 2.2500 4.1750 2.1400 4.1300 2.1400
                 4.1300 2.1300 3.0700 2.1300 3.0700 2.0650 2.2750 2.0650 2.2750 1.6300 2.4250 1.6300
                 2.4250 0.8700 2.2750 0.8700 2.2750 0.6300 2.3950 0.6300 2.3950 0.7500 2.5450 0.7500
                 2.5450 1.7500 2.3950 1.7500 2.3950 1.9450 3.1900 1.9450 3.1900 2.0100 4.2950 2.0100
                 4.2950 2.0200 5.0450 2.0200 5.0450 2.1200 5.8950 2.1200 5.8950 2.0200 6.6150 2.0200
                 6.6150 2.0700 6.7350 2.0700 ;
        POLYGON  6.1650 0.4800 6.0450 0.4800 6.0450 1.2800 5.5650 1.2800 5.5650 1.4000 5.4450 1.4000
                 5.4450 1.1600 5.9250 1.1600 5.9250 0.3600 6.1650 0.3600 ;
        POLYGON  5.8050 1.0400 5.3250 1.0400 5.3250 1.5200 5.5350 1.5200 5.5350 1.7600 5.4150 1.7600
                 5.4150 1.6400 5.2050 1.6400 5.2050 1.2800 3.4850 1.2800 3.4850 0.8200 3.0250 0.8200
                 3.0250 1.2200 2.9050 1.2200 2.9050 0.7000 3.6050 0.7000 3.6050 1.1600 5.2050 1.1600
                 5.2050 0.9200 5.6850 0.9200 5.6850 0.6200 5.8050 0.6200 ;
        POLYGON  5.4450 0.8000 5.0850 0.8000 5.0850 1.0400 4.2450 1.0400 4.2450 0.6200 4.3650 0.6200
                 4.3650 0.9200 4.9650 0.9200 4.9650 0.6800 5.4450 0.6800 ;
        POLYGON  5.0850 1.6600 4.8450 1.6600 4.8450 1.6500 3.6150 1.6500 3.6150 1.5300 4.9650 1.5300
                 4.9650 1.5400 5.0850 1.5400 ;
        POLYGON  4.8450 0.8000 4.6050 0.8000 4.6050 0.5000 4.1250 0.5000 4.1250 0.7200 3.9650 0.7200
                 3.9650 0.8000 3.7250 0.8000 3.7250 0.6800 3.8450 0.6800 3.8450 0.6000 4.0050 0.6000
                 4.0050 0.3800 4.7250 0.3800 4.7250 0.6800 4.8450 0.6800 ;
        POLYGON  3.8850 0.4800 3.7250 0.4800 3.7250 0.5600 2.7850 0.5600 2.7850 1.3400 2.8350 1.3400
                 2.8350 1.7200 2.7150 1.7200 2.7150 1.4600 2.6650 1.4600 2.6650 0.5600 2.5650 0.5600
                 2.5650 0.5100 2.1550 0.5100 2.1550 1.1100 1.8150 1.1100 1.8150 1.1500 1.5750 1.1500
                 1.5750 0.9900 2.0350 0.9900 2.0350 0.3900 2.6850 0.3900 2.6850 0.4400 3.6050 0.4400
                 3.6050 0.3600 3.8850 0.3600 ;
        POLYGON  1.1050 1.5800 0.9850 1.5800 0.9850 1.2000 0.3850 1.2000 0.3850 1.0800 0.9850 1.0800
                 0.9850 0.6800 1.1050 0.6800 ;
    END
END SDFFNSRXL

MACRO SDFFNSRX4
    CLASS CORE ;
    FOREIGN SDFFNSRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 16.2400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6750 0.3600 1.7950 1.4100 ;
        RECT  1.0150 0.3600 1.7950 0.4800 ;
        RECT  1.0150 0.9600 1.2350 1.2000 ;
        RECT  0.3750 0.9350 1.1350 1.0550 ;
        RECT  1.0150 0.3600 1.1350 1.2000 ;
        RECT  0.9400 0.5950 1.1350 1.0550 ;
        RECT  0.3750 0.9350 0.4950 1.1750 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.8950 1.4850 ;
        RECT  0.6500 1.1750 0.8000 1.4900 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1450 2.2500 1.4350 ;
        RECT  1.9950 0.9900 2.1150 1.2650 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0950 2.5400 1.4700 ;
        RECT  2.3900 0.9600 2.5100 1.4700 ;
        END
    END CKN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1550 0.9700 6.2750 1.2100 ;
        RECT  5.8150 0.9700 6.2750 1.0900 ;
        RECT  5.8150 0.9400 6.0750 1.0900 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5350 1.0900 7.4150 1.2100 ;
        RECT  6.3950 0.9400 6.6550 1.0900 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.8350 0.7400 13.0350 0.8600 ;
        RECT  12.7350 1.4200 12.8550 2.1900 ;
        RECT  12.5550 1.4200 12.8550 1.5400 ;
        RECT  11.9600 1.3000 12.6750 1.4200 ;
        RECT  11.9600 1.1750 12.1100 1.4350 ;
        RECT  11.9600 0.7400 12.0800 1.5400 ;
        RECT  11.8950 1.4200 12.0150 2.1900 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.7550 0.7400 14.9550 0.8600 ;
        RECT  14.4150 1.4200 14.5350 2.1900 ;
        RECT  14.2350 1.4200 14.5350 1.5400 ;
        RECT  13.7000 1.3000 14.3550 1.4200 ;
        RECT  13.5750 1.4200 13.8750 1.5400 ;
        RECT  13.7550 0.7400 13.8750 1.5400 ;
        RECT  13.7000 1.1750 13.8750 1.5400 ;
        RECT  13.5750 1.4200 13.6950 2.1900 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 16.2400 0.1800 ;
        RECT  15.3150 -0.1800 15.4350 0.7300 ;
        RECT  14.2350 -0.1800 14.4750 0.3800 ;
        RECT  13.2750 -0.1800 13.5150 0.3800 ;
        RECT  12.3150 -0.1800 12.5550 0.3800 ;
        RECT  11.3550 -0.1800 11.4750 0.8200 ;
        RECT  10.5150 -0.1800 10.6350 0.8600 ;
        RECT  7.0150 0.6100 7.2550 0.7300 ;
        RECT  7.1350 -0.1800 7.2550 0.7300 ;
        RECT  4.2200 -0.1800 4.4600 0.3200 ;
        RECT  1.9150 -0.1800 2.0350 0.8400 ;
        RECT  0.5550 -0.1800 0.6750 0.8150 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 16.2400 2.7900 ;
        RECT  14.8350 1.5400 14.9550 2.7900 ;
        RECT  13.9950 1.5400 14.1150 2.7900 ;
        RECT  13.1550 1.5400 13.2750 2.7900 ;
        RECT  12.3150 1.5400 12.4350 2.7900 ;
        RECT  11.4750 1.6400 11.5950 2.7900 ;
        RECT  10.6350 1.7000 10.7550 2.7900 ;
        RECT  9.5150 1.8800 9.7550 2.0000 ;
        RECT  9.5150 1.8800 9.6350 2.7900 ;
        RECT  6.3750 2.1300 6.6150 2.2500 ;
        RECT  6.3750 2.1300 6.4950 2.7900 ;
        RECT  4.8350 2.2000 5.0750 2.7900 ;
        RECT  4.2200 2.1700 4.3400 2.7900 ;
        RECT  4.1000 2.1700 4.3400 2.2900 ;
        RECT  2.1450 2.2300 2.2650 2.7900 ;
        RECT  0.6750 1.8500 0.7950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  15.8550 0.9200 15.6950 0.9200 15.6950 1.4200 15.3750 1.4200 15.3750 2.1900
                 15.2550 2.1900 15.2550 1.4200 14.6550 1.4200 14.6550 1.2800 14.8950 1.2800
                 14.8950 1.3000 15.5750 1.3000 15.5750 0.8000 15.7350 0.8000 15.7350 0.6800
                 15.8550 0.6800 ;
        POLYGON  15.4550 1.1800 15.2150 1.1800 15.2150 0.9700 15.0750 0.9700 15.0750 0.6200
                 11.7150 0.6200 11.7150 1.0600 11.2150 1.0600 11.2150 1.2800 11.7750 1.2800
                 11.7750 1.4000 11.2150 1.4000 11.2150 1.7600 11.1750 1.7600 11.1750 2.1600
                 11.0550 2.1600 11.0550 1.6400 11.0950 1.6400 11.0950 1.2400 9.9750 1.2400
                 9.9750 1.1200 10.9350 1.1200 10.9350 0.6800 11.0550 0.6800 11.0550 0.9400
                 11.5950 0.9400 11.5950 0.5000 15.1950 0.5000 15.1950 0.8500 15.3350 0.8500
                 15.3350 1.0600 15.4550 1.0600 ;
        POLYGON  10.9750 1.5200 8.5050 1.5200 8.5050 1.7700 8.3850 1.7700 8.3850 0.8700 8.3650 0.8700
                 8.3650 0.6300 8.4850 0.6300 8.4850 0.7500 8.5050 0.7500 8.5050 1.4000 10.7350 1.4000
                 10.7350 1.3600 10.9750 1.3600 ;
        POLYGON  10.3950 1.8800 9.8750 1.8800 9.8750 1.7600 8.7450 1.7600 8.7450 1.6400 9.9950 1.6400
                 9.9950 1.7600 10.3950 1.7600 ;
        POLYGON  10.2150 0.8600 10.0950 0.8600 10.0950 0.5600 9.4350 0.5600 9.4350 0.8000 9.1950 0.8000
                 9.1950 0.6800 9.3150 0.6800 9.3150 0.4400 10.2150 0.4400 ;
        POLYGON  9.8550 0.8000 9.6750 0.8000 9.6750 1.0400 8.8650 1.0400 8.8650 0.6300 8.9850 0.6300
                 8.9850 0.9200 9.5550 0.9200 9.5550 0.6800 9.8550 0.6800 ;
        POLYGON  9.5950 1.2800 8.6250 1.2800 8.6250 0.5100 7.6850 0.5100 7.6850 0.7400 7.6750 0.7400
                 7.6750 1.4100 7.6950 1.4100 7.6950 1.5300 7.4550 1.5300 7.4550 1.4100 7.5550 1.4100
                 7.5550 0.9700 6.7750 0.9700 6.7750 0.4800 6.1950 0.4800 6.1950 0.3600 6.8950 0.3600
                 6.8950 0.8500 7.3750 0.8500 7.3750 0.6200 7.5650 0.6200 7.5650 0.3900 8.7450 0.3900
                 8.7450 1.1600 9.5950 1.1600 ;
        POLYGON  9.3250 2.0500 9.0850 2.0500 9.0850 2.0100 6.9750 2.0100 6.9750 1.7700 5.6750 1.7700
                 5.6750 1.5700 4.9800 1.5700 4.9800 1.3300 5.1000 1.3300 5.1000 1.4500 5.7950 1.4500
                 5.7950 1.6500 7.0950 1.6500 7.0950 1.8900 8.1450 1.8900 8.1450 1.2300 8.0850 1.2300
                 8.0850 0.9900 8.2050 0.9900 8.2050 1.1100 8.2650 1.1100 8.2650 1.8900 9.2050 1.8900
                 9.2050 1.9300 9.3250 1.9300 ;
        POLYGON  8.3050 2.2500 6.7350 2.2500 6.7350 2.0100 5.4350 2.0100 5.4350 1.8100 4.5800 1.8100
                 4.5800 1.6900 4.7000 1.6900 4.7000 1.4400 3.7400 1.4400 3.7400 1.5600 3.6200 1.5600
                 3.6200 1.3200 4.7150 1.3200 4.7150 0.8400 4.6350 0.8400 4.6350 0.7200 4.8750 0.7200
                 4.8750 0.8400 4.8350 0.8400 4.8350 1.4400 4.8200 1.4400 4.8200 1.6900 5.5550 1.6900
                 5.5550 1.8900 6.8550 1.8900 6.8550 2.1300 8.3050 2.1300 ;
        POLYGON  8.0650 0.8700 7.9650 0.8700 7.9650 1.5300 8.0250 1.5300 8.0250 1.7700 7.2150 1.7700
                 7.2150 1.5300 5.9150 1.5300 5.9150 1.3300 5.5750 1.3300 5.5750 1.1000 4.9950 1.1000
                 4.9950 0.5600 3.9800 0.5600 3.9800 0.4800 3.8600 0.4800 3.8600 0.3600 4.1000 0.3600
                 4.1000 0.4400 5.1150 0.4400 5.1150 0.9800 5.5750 0.9800 5.5750 0.6800 5.8350 0.6800
                 5.8350 0.8000 5.6950 0.8000 5.6950 1.2100 6.0350 1.2100 6.0350 1.4100 7.3350 1.4100
                 7.3350 1.6500 7.8450 1.6500 7.8450 0.7500 7.9450 0.7500 7.9450 0.6300 8.0650 0.6300 ;
        POLYGON  6.2550 0.8000 5.9550 0.8000 5.9550 0.5600 5.4550 0.5600 5.4550 0.6200 5.3550 0.6200
                 5.3550 0.8600 5.2350 0.8600 5.2350 0.5000 5.3350 0.5000 5.3350 0.4400 6.0750 0.4400
                 6.0750 0.6800 6.2550 0.6800 ;
        POLYGON  5.9200 2.2500 5.1950 2.2500 5.1950 2.0500 3.4000 2.0500 3.4000 1.8000 3.3800 1.8000
                 3.3800 0.6200 3.5000 0.6200 3.5000 1.6800 3.5200 1.6800 3.5200 1.9300 5.3150 1.9300
                 5.3150 2.1300 5.9200 2.1300 ;
        POLYGON  4.5950 1.1600 3.8000 1.1600 3.8000 1.2000 3.6800 1.2000 3.6800 1.1600 3.6200 1.1600
                 3.6200 0.5000 3.2600 0.5000 3.2600 1.5600 3.1400 1.5600 3.1400 0.5000 2.5950 0.5000
                 2.5950 0.7200 2.7800 0.7200 2.7800 1.7100 2.7100 1.7100 2.7100 1.8300 2.5900 1.8300
                 2.5900 1.5900 2.6600 1.5900 2.6600 0.8400 2.4750 0.8400 2.4750 0.3800 3.7400 0.3800
                 3.7400 0.9600 3.8000 0.9600 3.8000 1.0400 4.5950 1.0400 ;
        POLYGON  3.1000 2.0700 1.4150 2.0700 1.4150 0.8400 1.2550 0.8400 1.2550 0.6000 1.3750 0.6000
                 1.3750 0.7200 1.5350 0.7200 1.5350 1.9500 2.9800 1.9500 2.9800 1.8300 2.9000 1.8300
                 2.9000 0.6200 3.0200 0.6200 3.0200 1.7100 3.1000 1.7100 ;
        POLYGON  1.2950 1.7300 0.3750 1.7300 0.3750 1.9700 0.2550 1.9700 0.2550 1.8500 0.1350 1.8500
                 0.1350 0.5750 0.2550 0.5750 0.2550 1.6100 1.1750 1.6100 1.1750 1.4100 1.2950 1.4100 ;
    END
END SDFFNSRX4

MACRO SDFFNSRX2
    CLASS CORE ;
    FOREIGN SDFFNSRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.5000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.1650 2.5950 1.3800 ;
        RECT  2.3350 0.9750 2.4550 1.3800 ;
        END
    END CKN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6700 1.3300 11.8200 1.7250 ;
        RECT  11.7000 1.0450 11.8200 1.7250 ;
        END
    END RN
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0800 0.8700 1.4350 ;
        RECT  0.7500 1.0750 0.8700 1.4350 ;
        END
    END SI
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.9750 1.9600 1.4450 ;
        RECT  1.8100 0.9750 1.9300 1.6150 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.7668  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 6.3900  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2900 0.9900 5.6700 1.1200 ;
        RECT  5.2900 0.8850 5.4400 1.1700 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0900 0.7550 1.2100 0.9950 ;
        RECT  0.9400 0.5950 1.0900 0.9550 ;
        RECT  0.3700 0.8350 1.2100 0.9550 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.4000 0.6800 12.5200 2.2050 ;
        RECT  12.2500 1.4650 12.5200 1.7250 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.2400 1.5450 13.4800 1.6650 ;
        RECT  13.3000 0.6800 13.4200 1.0850 ;
        RECT  13.2400 0.9650 13.3600 1.6650 ;
        RECT  13.0650 1.2300 13.3600 1.3800 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.5000 0.1800 ;
        RECT  13.7200 -0.1800 13.8400 0.9200 ;
        RECT  12.8800 -0.1800 13.0000 0.7300 ;
        RECT  11.8600 -0.1800 12.1000 0.3200 ;
        RECT  10.7500 -0.1800 10.8700 0.7800 ;
        RECT  6.0300 -0.1800 6.1500 0.8600 ;
        RECT  3.2500 -0.1800 3.4900 0.7400 ;
        RECT  2.0500 0.4950 2.2900 0.6150 ;
        RECT  2.1700 -0.1800 2.2900 0.6150 ;
        RECT  0.5900 -0.1800 0.7100 0.6750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.5000 2.7900 ;
        RECT  13.7200 2.0250 13.9600 2.1450 ;
        RECT  13.7200 2.0250 13.8400 2.7900 ;
        RECT  12.7600 2.0250 13.0000 2.1450 ;
        RECT  12.7600 2.0250 12.8800 2.7900 ;
        RECT  11.9800 1.8450 12.1000 2.7900 ;
        RECT  10.8100 2.2000 10.9300 2.7900 ;
        RECT  9.2900 1.9400 9.4100 2.7900 ;
        RECT  6.8900 1.9800 7.1300 2.1300 ;
        RECT  6.8900 1.9800 7.0100 2.7900 ;
        RECT  5.5700 1.8000 5.6900 2.7900 ;
        RECT  3.3000 1.7200 3.5400 1.8400 ;
        RECT  3.3000 1.7200 3.4200 2.7900 ;
        RECT  1.8700 1.7350 1.9900 2.7900 ;
        RECT  0.5300 2.2300 0.6500 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.3200 2.0850 14.2000 2.0850 14.2000 1.3250 13.5000 1.3250 13.5000 1.2050
                 14.1400 1.2050 14.1400 0.6800 14.2600 0.6800 14.2600 1.2050 14.3200 1.2050 ;
        POLYGON  14.0800 1.9050 12.8250 1.9050 12.8250 1.4550 12.6400 1.4550 12.6400 0.5600
                 12.2800 0.5600 12.2800 1.2600 12.1600 1.2600 12.1600 0.5600 11.2900 0.5600
                 11.2900 0.6800 11.3100 0.6800 11.3100 1.5200 11.2900 1.5200 11.2900 1.8400
                 11.1700 1.8400 11.1700 1.4000 11.1900 1.4000 11.1900 1.0200 10.2100 1.0200
                 10.2100 1.1000 10.0900 1.1000 10.0900 0.8600 10.2100 0.8600 10.2100 0.9000
                 11.1700 0.9000 11.1700 0.4400 12.7600 0.4400 12.7600 1.2150 12.9450 1.2150
                 12.9450 1.7850 13.9600 1.7850 13.9600 1.5050 14.0800 1.5050 ;
        POLYGON  11.6800 0.9250 11.5500 0.9250 11.5500 1.8450 11.6800 1.8450 11.6800 2.0850
                 11.5600 2.0850 11.5600 2.0800 10.7900 2.0800 10.7900 1.8200 10.1150 1.8200
                 10.1150 2.0100 9.7700 2.0100 9.7700 1.8900 9.9950 1.8900 9.9950 1.7000 10.9100 1.7000
                 10.9100 1.9600 11.4300 1.9600 11.4300 0.8050 11.5600 0.8050 11.5600 0.6800
                 11.6800 0.6800 ;
        POLYGON  11.0700 1.2600 10.9500 1.2600 10.9500 1.3400 8.4500 1.3400 8.4500 1.7200 8.3300 1.7200
                 8.3300 0.6800 8.5700 0.6800 8.5700 0.8000 8.4500 0.8000 8.4500 1.2200 10.8300 1.2200
                 10.8300 1.1400 11.0700 1.1400 ;
        POLYGON  10.6700 2.0600 10.5500 2.0600 10.5500 2.2500 9.5300 2.2500 9.5300 1.8200 9.1700 1.8200
                 9.1700 1.9000 8.9050 1.9000 8.9050 1.9600 8.4500 1.9600 8.4500 2.1400 7.2500 2.1400
                 7.2500 1.8600 6.7700 1.8600 6.7700 2.2500 5.8900 2.2500 5.8900 2.1300 6.6500 2.1300
                 6.6500 1.7400 7.3700 1.7400 7.3700 2.0200 8.3300 2.0200 8.3300 1.8400 8.7850 1.8400
                 8.7850 1.7800 9.0500 1.7800 9.0500 1.7000 9.6500 1.7000 9.6500 2.1300 10.4300 2.1300
                 10.4300 1.9400 10.6700 1.9400 ;
        POLYGON  10.5100 1.5800 8.9300 1.5800 8.9300 1.6600 8.6900 1.6600 8.6900 1.5400 8.8100 1.5400
                 8.8100 1.4600 10.5100 1.4600 ;
        POLYGON  10.4500 0.7800 10.3300 0.7800 10.3300 0.5400 10.2100 0.5400 10.2100 0.4800
                 9.7300 0.4800 9.7300 0.5400 9.6100 0.5400 9.6100 0.7800 9.4900 0.7800 9.4900 0.4200
                 9.6100 0.4200 9.6100 0.3600 10.3300 0.3600 10.3300 0.4200 10.4500 0.4200 ;
        POLYGON  10.0900 0.7200 9.9700 0.7200 9.9700 1.0200 8.8100 1.0200 8.8100 0.6200 8.9300 0.6200
                 8.9300 0.9000 9.8500 0.9000 9.8500 0.6000 10.0900 0.6000 ;
        POLYGON  8.7100 0.4800 8.2100 0.4800 8.2100 1.9000 7.4900 1.9000 7.4900 1.6200 6.5300 1.6200
                 6.5300 2.0100 5.8100 2.0100 5.8100 1.6800 5.2400 1.6800 5.2400 2.0000 5.0900 2.0000
                 5.0900 2.2000 4.8500 2.2000 4.8500 2.0000 3.7800 2.0000 3.7800 1.6400 3.8700 1.6400
                 3.8700 0.8600 3.8500 0.8600 3.8500 0.7400 4.0900 0.7400 4.0900 0.8600 3.9900 0.8600
                 3.9900 1.7600 3.9000 1.7600 3.9000 1.8800 4.4700 1.8800 4.4700 1.4000 4.4900 1.4000
                 4.4900 0.9800 4.6100 0.9800 4.6100 1.5200 4.5900 1.5200 4.5900 1.8800 5.1200 1.8800
                 5.1200 1.5600 5.9300 1.5600 5.9300 1.8900 6.4100 1.8900 6.4100 1.5000 7.6100 1.5000
                 7.6100 1.7800 8.0900 1.7800 8.0900 0.3600 8.7100 0.3600 ;
        POLYGON  7.9700 1.6600 7.7300 1.6600 7.7300 1.5400 7.8500 1.5400 7.8500 1.3800 6.1700 1.3800
                 6.1700 1.6500 6.2900 1.6500 6.2900 1.7700 6.0500 1.7700 6.0500 1.4400 5.2100 1.4400
                 5.2100 1.3200 6.0500 1.3200 6.0500 1.2600 6.8700 1.2600 6.8700 0.6200 6.9900 0.6200
                 6.9900 1.2600 7.8500 1.2600 7.8500 0.6200 7.9700 0.6200 ;
        POLYGON  7.4100 0.8600 7.2900 0.8600 7.2900 0.5000 6.7500 0.5000 6.7500 0.6200 6.5700 0.6200
                 6.5700 0.8600 6.4500 0.8600 6.4500 0.5000 6.6300 0.5000 6.6300 0.3800 7.4100 0.3800 ;
        POLYGON  6.6900 1.1400 5.7900 1.1400 5.7900 0.7650 4.9500 0.7650 4.9500 1.7600 4.7100 1.7600
                 4.7100 1.6400 4.8300 1.6400 4.8300 0.8000 4.7100 0.8000 4.7100 0.6800 4.8300 0.6800
                 4.8300 0.6450 5.9100 0.6450 5.9100 1.0200 6.6900 1.0200 ;
        POLYGON  4.4500 0.8600 4.3500 0.8600 4.3500 1.7600 4.1100 1.7600 4.1100 1.6400 4.2300 1.6400
                 4.2300 0.7400 4.3300 0.7400 4.3300 0.6200 3.7300 0.6200 3.7300 0.9800 3.0100 0.9800
                 3.0100 0.4950 2.5300 0.4950 2.5300 0.8550 1.8100 0.8550 1.8100 0.6350 1.4500 0.6350
                 1.4500 1.9150 1.1700 1.9150 1.1700 1.7950 1.3300 1.7950 1.3300 0.4350 1.4500 0.4350
                 1.4500 0.5150 1.9300 0.5150 1.9300 0.7350 2.4100 0.7350 2.4100 0.3750 3.1300 0.3750
                 3.1300 0.8600 3.6100 0.8600 3.6100 0.5000 4.4500 0.5000 ;
        POLYGON  3.7500 1.2200 2.8900 1.2200 2.8900 1.7950 2.2300 1.7950 2.2300 1.6750 2.7700 1.6750
                 2.7700 0.7350 2.6500 0.7350 2.6500 0.6150 2.8900 0.6150 2.8900 1.1000 3.7500 1.1000 ;
        POLYGON  1.6900 2.1550 0.9300 2.1550 0.9300 1.6750 0.2550 1.6750 0.2550 1.8300 0.1350 1.8300
                 0.1350 1.7100 0.1300 1.7100 0.1300 0.5950 0.1700 0.5950 0.1700 0.4350 0.2900 0.4350
                 0.2900 0.7150 0.2500 0.7150 0.2500 1.5550 1.0900 1.5550 1.0900 1.2950 1.2100 1.2950
                 1.2100 1.6750 1.0500 1.6750 1.0500 2.0350 1.5700 2.0350 1.5700 0.7550 1.6900 0.7550 ;
    END
END SDFFNSRX2

MACRO SDFFNSRX1
    CLASS CORE ;
    FOREIGN SDFFNSRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.0500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9050 1.2100 2.1450 1.3850 ;
        RECT  1.7550 1.2300 2.0150 1.4300 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7350 2.1300 7.5750 2.2500 ;
        RECT  6.7350 1.8000 6.8550 2.2500 ;
        RECT  5.1050 1.8000 6.8550 1.9200 ;
        RECT  5.1050 1.4000 5.2250 1.9200 ;
        RECT  3.6350 1.4000 5.2250 1.5200 ;
        RECT  3.6350 1.2300 3.7550 1.5200 ;
        RECT  3.3350 1.2700 3.7550 1.3900 ;
        RECT  3.4950 1.2300 3.7550 1.3900 ;
        END
    END SN
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5600 1.0300 10.6800 1.4650 ;
        RECT  10.5100 1.0300 10.6800 1.4450 ;
        END
    END CKN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.8000 1.4650 11.0250 1.7700 ;
        RECT  10.8300 1.4550 11.0250 1.7700 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.1950 1.4000 12.4550 1.6700 ;
        RECT  12.1900 1.4000 12.4550 1.6500 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.9500 1.1600 12.7500 1.2800 ;
        RECT  12.1950 0.9400 12.4550 1.2800 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 1.2950 1.4850 2.1400 ;
        RECT  1.3650 0.6100 1.4850 0.8500 ;
        RECT  1.2300 1.1750 1.4250 1.4350 ;
        RECT  1.3050 0.7300 1.4250 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.0500 0.1800 ;
        RECT  12.1900 -0.1800 12.3100 0.7300 ;
        RECT  10.8500 0.5500 11.0900 0.6700 ;
        RECT  10.9700 -0.1800 11.0900 0.6700 ;
        RECT  9.6500 -0.1800 9.8900 0.3400 ;
        RECT  7.8150 -0.1800 7.9350 0.8600 ;
        RECT  3.0150 -0.1800 3.1350 0.3800 ;
        RECT  1.7850 -0.1800 1.9050 0.8500 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.0500 2.7900 ;
        RECT  12.3050 2.0300 12.5450 2.1500 ;
        RECT  12.3050 2.0300 12.4250 2.7900 ;
        RECT  10.8650 1.9500 10.9850 2.7900 ;
        RECT  9.8850 1.6000 10.0050 2.7900 ;
        RECT  7.6950 2.1300 7.9350 2.2500 ;
        RECT  7.6950 2.1300 7.8150 2.7900 ;
        RECT  6.0350 2.2900 6.2750 2.7900 ;
        RECT  4.3550 2.1200 4.5950 2.2400 ;
        RECT  4.3550 2.1200 4.4750 2.7900 ;
        RECT  3.0750 1.7500 3.1950 2.7900 ;
        RECT  1.7850 1.5500 1.9050 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.9900 1.9700 12.9050 1.9700 12.9050 2.0900 12.7850 2.0900 12.7850 1.9100
                 11.9250 1.9100 11.9250 2.2500 11.1450 2.2500 11.1450 1.0300 11.5900 1.0300
                 11.5900 1.1500 11.2650 1.1500 11.2650 2.1300 11.8050 2.1300 11.8050 1.5100
                 11.9250 1.5100 11.9250 1.7900 12.8700 1.7900 12.8700 0.7300 12.7300 0.7300
                 12.7300 0.4900 12.8500 0.4900 12.8500 0.6100 12.9900 0.6100 ;
        POLYGON  11.8300 1.3900 11.6850 1.3900 11.6850 2.0100 11.4450 2.0100 11.4450 1.2700
                 11.7100 1.2700 11.7100 0.7300 11.4050 0.7300 11.4050 0.9100 10.6100 0.9100
                 10.6100 0.4800 10.1300 0.4800 10.1300 0.5800 9.6000 0.5800 9.6000 0.6200 8.9950 0.6200
                 8.9950 0.7400 9.2750 0.7400 9.2750 1.8900 9.1950 1.8900 9.1950 2.0100 9.0750 2.0100
                 9.0750 1.7700 9.1550 1.7700 9.1550 0.8600 8.8750 0.8600 8.8750 0.5000 9.4800 0.5000
                 9.4800 0.4600 10.0100 0.4600 10.0100 0.3600 10.7300 0.3600 10.7300 0.7900
                 11.2850 0.7900 11.2850 0.6100 11.5500 0.6100 11.5500 0.4900 11.6700 0.4900
                 11.6700 0.6100 11.8300 0.6100 ;
        POLYGON  10.4900 0.7200 10.3900 0.7200 10.3900 1.5650 10.4400 1.5650 10.4400 2.0700
                 10.3200 2.0700 10.3200 1.6850 10.2700 1.6850 10.2700 1.2200 9.8350 1.2200
                 9.8350 1.3400 9.7150 1.3400 9.7150 1.1000 10.2700 1.1000 10.2700 0.7200 10.2500 0.7200
                 10.2500 0.6000 10.4900 0.6000 ;
        POLYGON  9.6350 0.8600 9.5850 0.8600 9.5850 2.2500 8.8350 2.2500 8.8350 2.2200 8.2350 2.2200
                 8.2350 2.0100 6.9750 2.0100 6.9750 1.6800 6.7550 1.6800 6.7550 1.5600 6.3650 1.5600
                 6.3650 1.2300 6.4850 1.2300 6.4850 1.4400 6.8750 1.4400 6.8750 1.5600 7.0950 1.5600
                 7.0950 1.8900 8.2350 1.8900 8.2350 1.4800 8.4350 1.4800 8.4350 1.7200 8.3550 1.7200
                 8.3550 2.1000 8.8350 2.1000 8.8350 1.1200 8.7950 1.1200 8.7950 1.0000 9.0350 1.0000
                 9.0350 1.1200 8.9550 1.1200 8.9550 2.1300 9.4650 2.1300 9.4650 0.8600 9.3950 0.8600
                 9.3950 0.7400 9.6350 0.7400 ;
        POLYGON  8.7150 1.9800 8.4750 1.9800 8.4750 1.8600 8.5550 1.8600 8.5550 1.2000 7.2350 1.2000
                 7.2350 0.9600 7.3550 0.9600 7.3550 1.0800 8.5550 1.0800 8.5550 0.8600 8.4550 0.8600
                 8.4550 0.6200 8.5750 0.6200 8.5750 0.7400 8.6750 0.7400 8.6750 1.8600 8.7150 1.8600 ;
        POLYGON  8.1150 1.4400 7.3350 1.4400 7.3350 1.6500 7.4550 1.6500 7.4550 1.7700 7.2150 1.7700
                 7.2150 1.4400 6.9950 1.4400 6.9950 1.1100 6.2450 1.1100 6.2450 1.6400 5.7650 1.6400
                 5.7650 1.5200 6.1250 1.5200 6.1250 1.0200 5.8650 1.0200 5.8650 0.6200 5.9850 0.6200
                 5.9850 0.9000 6.2450 0.9000 6.2450 0.9900 6.9750 0.9900 6.9750 0.6200 7.0950 0.6200
                 7.0950 0.9900 7.1150 0.9900 7.1150 1.3200 8.1150 1.3200 ;
        POLYGON  7.5750 0.8000 7.3350 0.8000 7.3350 0.5000 6.8550 0.5000 6.8550 0.6800 6.7350 0.6800
                 6.7350 0.8000 6.4950 0.8000 6.4950 0.6800 6.6150 0.6800 6.6150 0.5600 6.7350 0.5600
                 6.7350 0.3800 7.4550 0.3800 7.4550 0.6800 7.5750 0.6800 ;
        POLYGON  6.6150 2.1700 4.7150 2.1700 4.7150 2.0000 4.2300 2.0000 4.2300 2.1300 4.2350 2.1300
                 4.2350 2.2500 3.9950 2.2500 3.9950 2.1200 3.3150 2.1200 3.3150 1.6300 2.9550 1.6300
                 2.9550 2.1100 2.2650 2.1100 2.2650 1.9100 2.2050 1.9100 2.2050 1.6700 2.2650 1.6700
                 2.2650 0.6100 2.3850 0.6100 2.3850 1.9900 2.8350 1.9900 2.8350 1.5100 3.4350 1.5100
                 3.4350 2.0000 4.1100 2.0000 4.1100 1.8800 4.8350 1.8800 4.8350 2.0500 6.6150 2.0500 ;
        POLYGON  6.0050 1.3800 5.8850 1.3800 5.8850 1.2600 5.6250 1.2600 5.6250 0.4800 5.1850 0.4800
                 5.1850 0.3600 5.7450 0.3600 5.7450 1.1400 6.0050 1.1400 ;
        POLYGON  5.5850 1.6400 5.3450 1.6400 5.3450 1.5200 5.3850 1.5200 5.3850 1.2800 3.9150 1.2800
                 3.9150 1.1100 3.0350 1.1100 3.0350 1.2400 2.9150 1.2400 2.9150 0.9900 4.0350 0.9900
                 4.0350 1.1600 5.3850 1.1600 5.3850 0.6200 5.5050 0.6200 5.5050 1.5200 5.5850 1.5200 ;
        POLYGON  5.0850 0.9200 4.9950 0.9200 4.9950 1.0400 4.1550 1.0400 4.1550 0.6200 4.2750 0.6200
                 4.2750 0.9200 4.8750 0.9200 4.8750 0.8000 4.9650 0.8000 4.9650 0.6200 5.0850 0.6200 ;
        POLYGON  4.9850 1.7600 3.6750 1.7600 3.6750 1.8800 3.5550 1.8800 3.5550 1.6400 4.9850 1.6400 ;
        POLYGON  4.7550 0.8000 4.5150 0.8000 4.5150 0.5000 4.0350 0.5000 4.0350 0.7200 3.7350 0.7200
                 3.7350 0.8000 3.4950 0.8000 3.4950 0.6800 3.6150 0.6800 3.6150 0.6000 3.9150 0.6000
                 3.9150 0.3800 4.6350 0.3800 4.6350 0.6800 4.7550 0.6800 ;
        POLYGON  3.7950 0.4800 3.3750 0.4800 3.3750 0.7500 3.1100 0.7500 3.1100 0.8700 2.7750 0.8700
                 2.7750 0.9000 2.7150 0.9000 2.7150 1.8700 2.5950 1.8700 2.5950 0.7500 2.6550 0.7500
                 2.6550 0.4900 2.1450 0.4900 2.1450 1.0900 1.7850 1.0900 1.7850 1.1100 1.5450 1.1100
                 1.5450 0.9700 2.0250 0.9700 2.0250 0.3700 2.7750 0.3700 2.7750 0.7500 2.9900 0.7500
                 2.9900 0.6300 3.2550 0.6300 3.2550 0.3600 3.7950 0.3600 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END SDFFNSRX1

MACRO SDFFHQX8
    CLASS CORE ;
    FOREIGN SDFFHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 1.3450 2.7750 2.1900 ;
        RECT  2.6550 0.6650 2.7750 0.9850 ;
        RECT  2.6350 0.8650 2.7550 1.4650 ;
        RECT  0.0700 1.0250 2.7550 1.1450 ;
        RECT  1.8150 0.6650 1.9350 2.1900 ;
        RECT  0.9750 0.6650 1.0950 2.1850 ;
        RECT  0.1350 0.6650 0.2550 2.1850 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 1.1550 5.2050 1.3800 ;
        RECT  5.0850 0.9800 5.2050 1.3800 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5350 1.2000 9.6550 1.4400 ;
        RECT  9.3500 1.2000 9.6550 1.4350 ;
        RECT  9.3500 1.1750 9.5000 1.4350 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7450 1.2100 11.1150 1.3950 ;
        RECT  10.7450 1.2100 11.0050 1.4200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.2750 0.9700 11.3950 1.2100 ;
        RECT  11.0350 0.9400 11.2950 1.0900 ;
        RECT  10.2750 0.9700 11.3950 1.0900 ;
        RECT  10.0150 1.0000 10.3950 1.1200 ;
        RECT  10.0150 1.0000 10.1350 1.4400 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  11.0750 -0.1800 11.1950 0.8200 ;
        RECT  9.7950 -0.1800 9.9150 0.6400 ;
        RECT  7.4250 -0.1800 7.6650 0.3700 ;
        RECT  5.3250 -0.1800 5.5650 0.3800 ;
        RECT  3.9150 -0.1800 4.0350 0.6500 ;
        RECT  3.0750 -0.1800 3.1950 0.6500 ;
        RECT  2.2350 -0.1800 2.3550 0.6550 ;
        RECT  1.3950 -0.1800 1.5150 0.6550 ;
        RECT  0.5550 -0.1800 0.6750 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  10.9150 1.7800 11.0350 2.7900 ;
        RECT  9.5350 1.8500 9.6550 2.7900 ;
        RECT  7.4250 2.0700 7.6650 2.1900 ;
        RECT  7.4250 2.0700 7.5450 2.7900 ;
        RECT  5.6450 2.1000 5.7650 2.7900 ;
        RECT  3.9750 1.5400 4.0950 2.7900 ;
        RECT  3.0750 1.4450 3.1950 2.7900 ;
        RECT  2.2350 1.4450 2.3550 2.7900 ;
        RECT  1.3950 1.4450 1.5150 2.7900 ;
        RECT  0.5550 1.4450 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6350 1.6800 11.5550 1.6800 11.5550 1.8000 11.4350 1.8000 11.4350 1.6600
                 10.4150 1.6600 10.4150 1.2400 10.5350 1.2400 10.5350 1.5400 11.5150 1.5400
                 11.5150 0.8500 11.4950 0.8500 11.4950 0.5800 11.6150 0.5800 11.6150 0.7300
                 11.6350 0.7300 ;
        POLYGON  10.5550 0.8500 10.1550 0.8500 10.1550 0.8800 9.8950 0.8800 9.8950 1.5600
                 10.2950 1.5600 10.2950 2.2100 10.1750 2.2100 10.1750 1.6800 8.9850 1.6800
                 8.9850 1.7600 8.7450 1.7600 8.7450 1.5300 8.8650 1.5300 8.8650 0.7200 8.7850 0.7200
                 8.7850 0.6000 9.0250 0.6000 9.0250 0.7200 8.9850 0.7200 8.9850 1.5600 9.7750 1.5600
                 9.7750 0.7600 10.0350 0.7600 10.0350 0.7300 10.4350 0.7300 10.4350 0.5900
                 10.5550 0.5900 ;
        POLYGON  9.4350 0.8300 9.3150 0.8300 9.3150 0.4800 8.6650 0.4800 8.6650 1.1500 8.7050 1.1500
                 8.7050 1.3900 8.6650 1.3900 8.6650 1.4100 8.6250 1.4100 8.6250 1.8800 9.1750 1.8800
                 9.1750 2.0300 9.2950 2.0300 9.2950 2.1500 9.0550 2.1500 9.0550 2.0000 8.5050 2.0000
                 8.5050 1.2900 8.5450 1.2900 8.5450 0.4800 8.0650 0.4800 8.0650 0.8800 8.1450 0.8800
                 8.1450 1.1200 7.9450 1.1200 7.9450 0.6100 7.1850 0.6100 7.1850 0.4800 6.7050 0.4800
                 6.7050 0.9700 6.9650 0.9700 6.9650 1.2100 6.8450 1.2100 6.8450 1.0900 6.5850 1.0900
                 6.5850 0.3600 7.3050 0.3600 7.3050 0.4900 7.9450 0.4900 7.9450 0.3600 9.4350 0.3600 ;
        POLYGON  8.4250 0.7200 8.3850 0.7200 8.3850 1.9900 8.2650 1.9900 8.2650 1.3600 7.4650 1.3600
                 7.4650 1.3100 7.3250 1.3100 7.3250 1.1900 7.5850 1.1900 7.5850 1.2400 8.2650 1.2400
                 8.2650 0.7200 8.1850 0.7200 8.1850 0.6000 8.4250 0.6000 ;
        POLYGON  8.2250 2.2500 7.9850 2.2500 7.9850 1.9500 7.0450 1.9500 7.0450 2.2300 5.9250 2.2300
                 5.9250 0.8600 4.8250 0.8600 4.8250 1.5000 5.2450 1.5000 5.2450 1.7400 5.1250 1.7400
                 5.1250 1.6200 4.7050 1.6200 4.7050 0.6000 4.9650 0.6000 4.9650 0.7400 6.0450 0.7400
                 6.0450 2.1100 6.5850 2.1100 6.5850 1.3300 6.4250 1.3300 6.4250 1.2100 6.7050 1.2100
                 6.7050 2.1100 6.9250 2.1100 6.9250 1.8300 8.1050 1.8300 8.1050 2.1300 8.2250 2.1300 ;
        POLYGON  7.8250 1.1200 7.7050 1.1200 7.7050 1.0700 7.2050 1.0700 7.2050 1.4500 7.1250 1.4500
                 7.1250 1.7100 7.0050 1.7100 7.0050 1.3300 7.0850 1.3300 7.0850 0.8500 6.8250 0.8500
                 6.8250 0.6000 7.0650 0.6000 7.0650 0.7300 7.2050 0.7300 7.2050 0.9500 7.7050 0.9500
                 7.7050 0.8800 7.8250 0.8800 ;
        POLYGON  6.4650 1.9900 6.3450 1.9900 6.3450 1.5700 6.1850 1.5700 6.1850 0.6200 5.0850 0.6200
                 5.0850 0.4800 4.2750 0.4800 4.2750 1.1800 4.1550 1.1800 4.1550 0.3600 5.2050 0.3600
                 5.2050 0.5000 6.3050 0.5000 6.3050 1.4500 6.4650 1.4500 ;
        POLYGON  5.7250 1.9800 4.5150 1.9800 4.5150 2.1900 4.3950 2.1900 4.3950 1.4200 3.6750 1.4200
                 3.6750 2.1900 3.5550 2.1900 3.5550 1.5400 3.4950 1.5400 3.4950 1.2250 2.8750 1.2250
                 2.8750 1.1050 3.4950 1.1050 3.4950 0.6000 3.6150 0.6000 3.6150 1.3000 4.3950 1.3000
                 4.3950 0.6000 4.5150 0.6000 4.5150 1.8600 5.6050 1.8600 5.6050 1.1300 5.7250 1.1300 ;
    END
END SDFFHQX8

MACRO SDFFHQX4
    CLASS CORE ;
    FOREIGN SDFFHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1850 0.6300 2.3050 0.8700 ;
        RECT  1.9650 1.3150 2.2050 1.6500 ;
        RECT  2.0850 0.7500 2.2050 1.6500 ;
        RECT  1.2300 1.3150 2.2050 1.4350 ;
        RECT  1.3450 0.6300 1.4650 0.8700 ;
        RECT  1.0050 1.5300 1.3800 1.6500 ;
        RECT  1.2300 1.1750 1.3800 1.6500 ;
        RECT  1.2600 0.7500 1.3800 1.6500 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1750 0.6850 1.2950 ;
        RECT  0.5650 1.0550 0.6850 1.2950 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5950 1.2000 7.7150 1.4400 ;
        RECT  7.3200 1.3150 7.7150 1.4350 ;
        RECT  7.3200 1.1750 7.4700 1.4350 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7150 1.2300 9.0600 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0050 0.9900 9.3750 1.1100 ;
        RECT  8.2350 0.9700 9.2650 1.0900 ;
        RECT  9.0050 0.9400 9.2650 1.1100 ;
        RECT  8.0750 1.1900 8.3550 1.3100 ;
        RECT  8.2350 0.9700 8.3550 1.3100 ;
        RECT  8.0750 1.1900 8.1950 1.4400 ;
        END
    END SE
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.1350 -0.1800 9.2550 0.8200 ;
        RECT  7.7550 -0.1800 7.8750 0.8300 ;
        RECT  5.4650 0.3900 5.7050 0.5100 ;
        RECT  5.5850 -0.1800 5.7050 0.5100 ;
        RECT  3.4450 -0.1800 3.5650 0.6800 ;
        RECT  2.6050 -0.1800 2.7250 0.6800 ;
        RECT  1.7650 -0.1800 1.8850 0.6800 ;
        RECT  0.9250 -0.1800 1.0450 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  8.9750 1.7950 9.0950 2.7900 ;
        RECT  7.5950 1.8500 7.7150 2.7900 ;
        RECT  5.4650 2.0700 5.7050 2.1900 ;
        RECT  5.4650 2.0700 5.5850 2.7900 ;
        RECT  3.4050 2.0100 3.6450 2.1300 ;
        RECT  3.4050 2.0100 3.5250 2.7900 ;
        RECT  2.4450 2.0100 2.6850 2.1300 ;
        RECT  2.4450 2.0100 2.5650 2.7900 ;
        RECT  1.4850 2.0100 1.7250 2.1300 ;
        RECT  1.4850 2.0100 1.6050 2.7900 ;
        RECT  0.5850 2.1100 0.7050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.6750 0.8200 9.6150 0.8200 9.6150 1.6800 9.5750 1.6800 9.5750 1.8000 9.4550 1.8000
                 9.4550 1.6750 8.4750 1.6750 8.4750 1.2400 8.5950 1.2400 8.5950 1.5550 9.4950 1.5550
                 9.4950 0.7000 9.5550 0.7000 9.5550 0.5800 9.6750 0.5800 ;
        POLYGON  8.6150 0.8500 8.1150 0.8500 8.1150 1.0700 7.9550 1.0700 7.9550 1.5600 8.3550 1.5600
                 8.3550 2.2100 8.2350 2.2100 8.2350 1.6800 7.0250 1.6800 7.0250 1.7600 6.7850 1.7600
                 6.7850 1.5300 6.9050 1.5300 6.9050 0.7200 6.8850 0.7200 6.8850 0.6000 7.1250 0.6000
                 7.1250 0.7200 7.0250 0.7200 7.0250 1.5600 7.8350 1.5600 7.8350 0.9500 7.9950 0.9500
                 7.9950 0.7300 8.4950 0.7300 8.4950 0.5900 8.6150 0.5900 ;
        POLYGON  7.4550 0.8300 7.3350 0.8300 7.3350 0.4800 6.7650 0.4800 6.7650 1.3900 6.6650 1.3900
                 6.6650 1.8800 7.2350 1.8800 7.2350 2.0300 7.3550 2.0300 7.3550 2.1500 7.1150 2.1500
                 7.1150 2.0000 6.5450 2.0000 6.5450 1.1500 6.6450 1.1500 6.6450 0.4800 6.1650 0.4800
                 6.1650 0.8800 6.1850 0.8800 6.1850 1.1200 6.0450 1.1200 6.0450 0.7500 5.2250 0.7500
                 5.2250 0.4800 4.7450 0.4800 4.7450 1.0000 4.6650 1.0000 4.6650 1.2500 4.1250 1.2500
                 4.1250 1.3700 4.0050 1.3700 4.0050 1.1300 4.5450 1.1300 4.5450 0.8800 4.6250 0.8800
                 4.6250 0.3600 5.3450 0.3600 5.3450 0.6300 6.0450 0.6300 6.0450 0.3600 7.4550 0.3600 ;
        POLYGON  6.5250 0.7200 6.4250 0.7200 6.4250 1.9900 6.3050 1.9900 6.3050 1.3600 5.4850 1.3600
                 5.4850 1.3100 5.3650 1.3100 5.3650 1.1900 5.6050 1.1900 5.6050 1.2400 6.3050 1.2400
                 6.3050 0.7200 6.2850 0.7200 6.2850 0.6000 6.5250 0.6000 ;
        POLYGON  6.2650 2.2500 6.0250 2.2500 6.0250 1.9500 4.9250 1.9500 4.9250 2.2300 3.8450 2.2300
                 3.8450 1.8900 0.1350 1.8900 0.1350 1.6750 0.1200 1.6750 0.1200 0.9350 0.3250 0.9350
                 0.3250 0.6300 0.4450 0.6300 0.4450 1.0550 0.2400 1.0550 0.2400 1.5550 0.2550 1.5550
                 0.2550 1.7700 3.9650 1.7700 3.9650 2.1100 4.8050 2.1100 4.8050 1.2300 4.8850 1.2300
                 4.8850 1.1100 5.0050 1.1100 5.0050 1.3500 4.9250 1.3500 4.9250 1.8300 6.1450 1.8300
                 6.1450 2.1300 6.2650 2.1300 ;
        POLYGON  5.9250 1.0700 5.2450 1.0700 5.2450 1.5900 5.1650 1.5900 5.1650 1.7100 5.0450 1.7100
                 5.0450 1.4700 5.1250 1.4700 5.1250 0.9900 4.8650 0.9900 4.8650 0.6000 5.1050 0.6000
                 5.1050 0.8700 5.2450 0.8700 5.2450 0.9500 5.9250 0.9500 ;
        POLYGON  4.5050 0.7200 3.8850 0.7200 3.8850 1.4900 4.2450 1.4900 4.2450 1.4700 4.3650 1.4700
                 4.3650 1.9900 4.2450 1.9900 4.2450 1.6100 3.7650 1.6100 3.7650 1.3700 3.1850 1.3700
                 3.1850 1.1300 3.3050 1.1300 3.3050 1.2500 3.7650 1.2500 3.7650 0.6000 4.5050 0.6000 ;
        POLYGON  3.6450 1.1300 3.5250 1.1300 3.5250 1.0100 3.0650 1.0100 3.0650 1.5300 3.1650 1.5300
                 3.1650 1.6500 2.9250 1.6500 2.9250 1.5300 2.9450 1.5300 2.9450 1.0100 2.5450 1.0100
                 2.5450 1.1900 2.4250 1.1900 2.4250 0.8900 2.9450 0.8900 2.9450 0.6600 3.0250 0.6600
                 3.0250 0.5400 3.1450 0.5400 3.1450 0.8900 3.6450 0.8900 ;
    END
END SDFFHQX4

MACRO SDFFHQX2
    CLASS CORE ;
    FOREIGN SDFFHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.4650 1.3350 1.5850 ;
        RECT  1.2150 1.3450 1.3350 1.5850 ;
        RECT  0.9400 1.4650 1.0900 1.7250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4850 0.9600 6.6800 1.2000 ;
        RECT  6.4500 0.8850 6.6750 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9000 1.0250 8.0600 1.4800 ;
        RECT  7.9400 1.0000 8.0600 1.4800 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4250 1.2300 8.6850 1.3800 ;
        RECT  8.4250 1.0700 8.5450 1.3800 ;
        RECT  8.3400 0.7600 8.4600 1.1900 ;
        RECT  8.2200 1.0700 8.5450 1.1900 ;
        RECT  7.3000 0.7600 8.4600 0.8800 ;
        RECT  7.5400 0.7600 7.7800 1.0900 ;
        RECT  7.0400 1.0000 7.4200 1.1200 ;
        RECT  7.3000 0.7600 7.4200 1.1200 ;
        RECT  7.0400 1.0000 7.1600 1.4400 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6800 0.6750 2.2050 ;
        RECT  0.3600 1.1750 0.6750 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.1000 -0.1800 8.2200 0.6400 ;
        RECT  6.8200 -0.1800 6.9400 0.6400 ;
        RECT  4.4300 0.3800 4.6700 0.5000 ;
        RECT  4.5500 -0.1800 4.6700 0.5000 ;
        RECT  2.5700 -0.1800 2.6900 0.6800 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  7.9400 1.8400 8.0600 2.7900 ;
        RECT  6.5600 1.5600 6.6800 2.7900 ;
        RECT  4.4300 2.0600 4.6700 2.1800 ;
        RECT  4.4300 2.0600 4.5500 2.7900 ;
        RECT  2.3100 2.0600 2.4300 2.7900 ;
        RECT  0.9750 1.8450 1.0950 2.7900 ;
        RECT  0.1350 1.5550 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.9250 1.7200 8.5400 1.7200 8.5400 1.8400 8.4200 1.8400 8.4200 1.7200 7.4400 1.7200
                 7.4400 1.2400 7.5600 1.2400 7.5600 1.6000 8.8050 1.6000 8.8050 0.9500 8.5800 0.9500
                 8.5800 0.5900 8.7000 0.5900 8.7000 0.8300 8.9250 0.8300 ;
        POLYGON  7.5800 0.6400 7.1800 0.6400 7.1800 0.8800 6.9200 0.8800 6.9200 1.5600 7.3200 1.5600
                 7.3200 2.2100 7.2000 2.2100 7.2000 1.6800 6.8000 1.6800 6.8000 1.4400 5.9900 1.4400
                 5.9900 1.5800 5.9500 1.5800 5.9500 1.7000 5.8300 1.7000 5.8300 1.4600 5.8700 1.4600
                 5.8700 0.7200 5.8300 0.7200 5.8300 0.6000 6.0700 0.6000 6.0700 0.7200 5.9900 0.7200
                 5.9900 1.3200 6.8000 1.3200 6.8000 0.7600 7.0600 0.7600 7.0600 0.5200 7.4600 0.5200
                 7.4600 0.4000 7.5800 0.4000 ;
        POLYGON  6.4600 0.6600 6.3400 0.6600 6.3400 0.4800 5.7100 0.4800 5.7100 1.1000 5.7500 1.1000
                 5.7500 1.3400 5.7100 1.3400 5.7100 1.9100 6.2600 1.9100 6.2600 2.0300 5.5900 2.0300
                 5.5900 0.4800 5.1100 0.4800 5.1100 0.9200 5.2300 0.9200 5.2300 1.0400 4.9900 1.0400
                 4.9900 0.7400 4.1900 0.7400 4.1900 0.4800 3.7100 0.4800 3.7100 0.9800 3.5700 0.9800
                 3.5700 1.2600 2.9900 1.2600 2.9900 1.3800 2.8700 1.3800 2.8700 1.1400 3.4500 1.1400
                 3.4500 0.8600 3.5900 0.8600 3.5900 0.3600 4.3100 0.3600 4.3100 0.6200 4.9900 0.6200
                 4.9900 0.3600 6.4600 0.3600 ;
        POLYGON  5.4700 1.9800 5.3500 1.9800 5.3500 1.3000 4.2900 1.3000 4.2900 1.1800 5.3500 1.1800
                 5.3500 0.7200 5.2300 0.7200 5.2300 0.6000 5.4700 0.6000 ;
        POLYGON  5.2500 2.2400 5.0100 2.2400 5.0100 1.9400 3.8900 1.9400 3.8900 2.2200 2.7100 2.2200
                 2.7100 1.9400 2.0350 1.9400 2.0350 1.9650 1.5150 1.9650 1.5150 2.0850 1.3950 2.0850
                 1.3950 1.8450 1.4550 1.8450 1.4550 0.6800 1.5750 0.6800 1.5750 1.8450 1.9150 1.8450
                 1.9150 1.8200 2.8300 1.8200 2.8300 2.1000 3.7700 2.1000 3.7700 1.2200 3.8100 1.2200
                 3.8100 1.1000 3.9300 1.1000 3.9300 1.3400 3.8900 1.3400 3.8900 1.8200 5.1300 1.8200
                 5.1300 2.1200 5.2500 2.1200 ;
        POLYGON  4.8700 1.0600 4.1700 1.0600 4.1700 1.5800 4.1300 1.5800 4.1300 1.7000 4.0100 1.7000
                 4.0100 1.4600 4.0500 1.4600 4.0500 0.9800 3.8300 0.9800 3.8300 0.6000 4.0700 0.6000
                 4.0700 0.8600 4.1700 0.8600 4.1700 0.9400 4.8700 0.9400 ;
        POLYGON  3.4700 0.7200 2.9300 0.7200 2.9300 1.0200 2.7500 1.0200 2.7500 1.5000 3.1100 1.5000
                 3.1100 1.4600 3.2300 1.4600 3.2300 1.9800 3.1100 1.9800 3.1100 1.6200 2.0700 1.6200
                 2.0700 1.3400 2.0500 1.3400 2.0500 1.1000 2.1900 1.1000 2.1900 1.5000 2.6300 1.5000
                 2.6300 0.9000 2.8100 0.9000 2.8100 0.6000 3.4700 0.6000 ;
        POLYGON  2.5100 1.3800 2.3900 1.3800 2.3900 0.9800 1.9300 0.9800 1.9300 1.4600 1.9500 1.4600
                 1.9500 1.7000 1.8300 1.7000 1.8300 1.5800 1.8100 1.5800 1.8100 0.5600 1.3350 0.5600
                 1.3350 1.1800 0.7950 1.1800 0.7950 1.0600 1.2150 1.0600 1.2150 0.4400 2.2700 0.4400
                 2.2700 0.8600 2.5100 0.8600 ;
    END
END SDFFHQX2

MACRO SDFFHQX1
    CLASS CORE ;
    FOREIGN SDFFHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7100 1.0900 0.8600 1.4250 ;
        RECT  0.6500 1.0950 0.8300 1.4350 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0650 0.9600 6.1850 1.2000 ;
        RECT  5.8700 0.9600 6.1850 1.1450 ;
        RECT  5.8700 0.8850 6.0200 1.1450 ;
        END
    END D
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.2100 7.6250 1.4100 ;
        RECT  7.2650 1.2100 7.5250 1.4350 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7650 0.9700 7.8850 1.2100 ;
        RECT  7.5550 0.9400 7.8150 1.0900 ;
        RECT  6.5450 0.9700 7.8850 1.0900 ;
        RECT  6.5450 0.9700 6.6650 1.4400 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.2950 0.2650 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.6650 -0.1800 7.7850 0.8200 ;
        RECT  6.0650 -0.1800 6.1850 0.6400 ;
        RECT  3.7950 0.3900 4.0350 0.5100 ;
        RECT  3.7950 -0.1800 3.9150 0.5100 ;
        RECT  2.0150 -0.1800 2.1350 0.6800 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.4450 1.7950 7.5650 2.7900 ;
        RECT  6.0650 1.5600 6.1850 2.7900 ;
        RECT  3.7950 2.0700 4.0350 2.1900 ;
        RECT  3.7950 2.0700 3.9150 2.7900 ;
        RECT  1.7150 2.0100 1.9550 2.1300 ;
        RECT  1.7150 2.0100 1.8350 2.7900 ;
        RECT  0.5650 1.8500 0.6850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2050 0.8200 8.1250 0.8200 8.1250 1.6800 8.0450 1.6800 8.0450 1.8000 7.9250 1.8000
                 7.9250 1.6750 6.9450 1.6750 6.9450 1.2400 7.0650 1.2400 7.0650 1.5550 8.0050 1.5550
                 8.0050 0.7000 8.0850 0.7000 8.0850 0.5800 8.2050 0.5800 ;
        POLYGON  7.1450 0.8500 6.4250 0.8500 6.4250 1.5600 6.8250 1.5600 6.8250 2.2100 6.7050 2.2100
                 6.7050 1.6800 6.3050 1.6800 6.3050 1.4400 5.3550 1.4400 5.3550 1.5900 5.2550 1.5900
                 5.2550 1.9900 5.1350 1.9900 5.1350 1.4700 5.2350 1.4700 5.2350 0.7200 5.1350 0.7200
                 5.1350 0.6000 5.3750 0.6000 5.3750 0.7200 5.3550 0.7200 5.3550 1.3200 6.3050 1.3200
                 6.3050 0.7300 7.0250 0.7300 7.0250 0.5900 7.1450 0.5900 ;
        POLYGON  5.7650 1.8600 5.6450 1.8600 5.6450 1.9800 5.4950 1.9800 5.4950 2.2300 4.8950 2.2300
                 4.8950 0.4800 4.4150 0.4800 4.4150 0.8400 4.5350 0.8400 4.5350 1.1000 4.4150 1.1000
                 4.4150 0.9600 4.2950 0.9600 4.2950 0.7500 3.5550 0.7500 3.5550 0.4800 3.0750 0.4800
                 3.0750 0.9800 3.0350 0.9800 3.0350 1.1000 3.0150 1.1000 3.0150 1.2700 2.4550 1.2700
                 2.4550 1.3900 2.3350 1.3900 2.3350 1.1500 2.8950 1.1500 2.8950 0.8600 2.9550 0.8600
                 2.9550 0.3600 3.6750 0.3600 3.6750 0.6300 4.2950 0.6300 4.2950 0.3600 5.7050 0.3600
                 5.7050 0.8100 5.5850 0.8100 5.5850 0.4800 5.0150 0.4800 5.0150 1.1100 5.1150 1.1100
                 5.1150 1.3500 5.0150 1.3500 5.0150 2.1100 5.3750 2.1100 5.3750 1.8600 5.5250 1.8600
                 5.5250 1.7400 5.7650 1.7400 ;
        POLYGON  4.7750 1.9900 4.6550 1.9900 4.6550 1.5600 3.7550 1.5600 3.7550 1.1300 3.8750 1.1300
                 3.8750 1.4400 4.6550 1.4400 4.6550 0.7200 4.5350 0.7200 4.5350 0.6000 4.7750 0.6000 ;
        POLYGON  4.5950 2.2500 4.3550 2.2500 4.3550 1.9500 3.2550 1.9500 3.2550 2.2300 2.0750 2.2300
                 2.0750 1.8900 1.1050 1.8900 1.1050 2.1000 0.9850 2.1000 0.9850 1.2900 1.0350 1.2900
                 1.0350 0.6800 1.1550 0.6800 1.1550 1.4100 1.1050 1.4100 1.1050 1.7700 2.1950 1.7700
                 2.1950 2.1100 3.1350 2.1100 3.1350 1.2300 3.2750 1.2300 3.2750 1.1100 3.3950 1.1100
                 3.3950 1.3500 3.2550 1.3500 3.2550 1.8300 4.4750 1.8300 4.4750 2.1300 4.5950 2.1300 ;
        POLYGON  4.1950 1.3200 4.0550 1.3200 4.0550 1.0100 3.6350 1.0100 3.6350 1.5900 3.4950 1.5900
                 3.4950 1.7100 3.3750 1.7100 3.3750 1.4700 3.5150 1.4700 3.5150 0.9900 3.1950 0.9900
                 3.1950 0.6000 3.4350 0.6000 3.4350 0.8700 3.6350 0.8700 3.6350 0.8900 4.1750 0.8900
                 4.1750 1.0800 4.1950 1.0800 ;
        POLYGON  2.8350 0.7200 2.3750 0.7200 2.3750 1.0300 2.2150 1.0300 2.2150 1.5100 2.5750 1.5100
                 2.5750 1.4700 2.6950 1.4700 2.6950 1.9900 2.5750 1.9900 2.5750 1.6300 1.5950 1.6300
                 1.5950 1.3700 1.5150 1.3700 1.5150 1.1300 1.7150 1.1300 1.7150 1.5100 2.0950 1.5100
                 2.0950 0.9100 2.2550 0.9100 2.2550 0.6000 2.8350 0.6000 ;
        POLYGON  1.9750 1.3900 1.8550 1.3900 1.8550 1.0100 1.3950 1.0100 1.3950 1.5300 1.4750 1.5300
                 1.4750 1.6500 1.2350 1.6500 1.2350 1.5300 1.2750 1.5300 1.2750 0.5600 0.9150 0.5600
                 0.9150 0.9700 0.5200 0.9700 0.5200 1.2400 0.4000 1.2400 0.4000 0.8500 0.7950 0.8500
                 0.7950 0.4400 1.7150 0.4400 1.7150 0.8900 1.9750 0.8900 ;
    END
END SDFFHQX1

MACRO OR4XL
    CLASS CORE ;
    FOREIGN OR4XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.0200 1.6750 1.4550 ;
        RECT  1.5350 1.0200 1.6600 1.4800 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1750 0.5100 1.6300 ;
        RECT  0.3600 1.1750 0.4800 1.6600 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1250 0.8200 1.5400 ;
        RECT  0.7000 1.1050 0.8200 1.5400 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0400 1.3300 1.1600 1.6600 ;
        RECT  0.9400 1.1750 1.0900 1.5100 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0550 2.4400 1.1750 ;
        RECT  2.3200 0.6600 2.4400 1.1750 ;
        RECT  2.1000 1.0550 2.2500 1.4350 ;
        RECT  2.1000 1.0550 2.2200 1.9600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.9000 -0.1800 2.0200 0.9000 ;
        RECT  1.0400 -0.1800 1.1600 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.6800 1.8400 1.8000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9800 1.7200 1.4000 1.7200 1.4000 1.9000 0.1600 1.9000 0.1600 1.7800 1.2800 1.7800
                 1.2800 0.9000 0.5600 0.9000 0.5600 0.6600 0.6800 0.6600 0.6800 0.7800 1.4800 0.7800
                 1.4800 0.6600 1.6000 0.6600 1.6000 0.9000 1.4000 0.9000 1.4000 1.6000 1.8600 1.6000
                 1.8600 1.3800 1.9800 1.3800 ;
    END
END OR4XL

MACRO OR4X8
    CLASS CORE ;
    FOREIGN OR4X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9500 2.1350 1.1300 ;
        RECT  1.7550 0.9400 2.0150 1.1300 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2550 1.2500 2.5950 1.3700 ;
        RECT  2.4750 0.9400 2.5950 1.3700 ;
        RECT  2.3350 0.9400 2.5950 1.0900 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.4900 2.9750 1.6100 ;
        RECT  2.8550 1.2400 2.9750 1.6100 ;
        RECT  0.6800 1.2800 1.0750 1.6100 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2050 1.5200 3.4650 1.6700 ;
        RECT  0.4100 1.7300 3.3350 1.8500 ;
        RECT  3.2150 1.2200 3.3350 1.8500 ;
        RECT  3.2050 1.5200 3.3350 1.8500 ;
        RECT  0.4100 1.2200 0.5300 1.8500 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3350 0.7150 6.6950 0.8350 ;
        RECT  6.4150 1.2300 6.5350 2.2100 ;
        RECT  4.0550 0.7650 6.4550 0.8850 ;
        RECT  5.6950 1.2300 6.5350 1.3500 ;
        RECT  5.6950 0.7650 6.0200 1.3500 ;
        RECT  3.8950 1.2750 5.8150 1.3950 ;
        RECT  5.6750 0.6450 5.7950 0.8850 ;
        RECT  5.5750 1.2750 5.6950 2.2100 ;
        RECT  4.7750 0.7150 5.0150 0.8850 ;
        RECT  4.7350 1.2750 4.8550 2.2100 ;
        RECT  3.9350 0.7150 4.1750 0.8350 ;
        RECT  3.8950 1.2750 4.0150 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  6.0950 -0.1800 6.2150 0.6450 ;
        RECT  5.2550 -0.1800 5.3750 0.6450 ;
        RECT  4.4150 -0.1800 4.5350 0.6450 ;
        RECT  3.5150 0.4600 3.7550 0.5800 ;
        RECT  3.5150 -0.1800 3.6350 0.5800 ;
        RECT  2.6750 0.4600 2.9150 0.5800 ;
        RECT  2.6750 -0.1800 2.7950 0.5800 ;
        RECT  1.8350 0.4600 2.0750 0.5800 ;
        RECT  1.8350 -0.1800 1.9550 0.5800 ;
        RECT  0.9950 0.4600 1.2350 0.5800 ;
        RECT  0.9950 -0.1800 1.1150 0.5800 ;
        RECT  0.2150 -0.1800 0.3350 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  5.9950 1.4700 6.1150 2.7900 ;
        RECT  5.1550 1.5150 5.2750 2.7900 ;
        RECT  4.3150 1.5150 4.4350 2.7900 ;
        RECT  3.3550 2.2100 3.5950 2.7900 ;
        RECT  0.4150 1.9700 0.5350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.5750 1.1550 3.7050 1.1550 3.7050 2.0900 2.1750 2.0900 2.1750 2.1500 1.9350 2.1500
                 1.9350 1.9700 3.5850 1.9700 3.5850 0.8200 0.6950 0.8200 0.6950 0.7700 0.5750 0.7700
                 0.5750 0.6500 0.8150 0.6500 0.8150 0.7000 1.4150 0.7000 1.4150 0.6500 1.6550 0.6500
                 1.6550 0.7000 2.2550 0.7000 2.2550 0.6500 2.4950 0.6500 2.4950 0.7000 3.0950 0.7000
                 3.0950 0.6500 3.3350 0.6500 3.3350 0.7000 3.7050 0.7000 3.7050 1.0350 5.5750 1.0350 ;
    END
END OR4X8

MACRO OR4X6
    CLASS CORE ;
    FOREIGN OR4X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9500 2.1350 1.1300 ;
        RECT  1.7550 0.9400 2.0150 1.1300 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2550 1.2500 2.5950 1.3700 ;
        RECT  2.4750 0.9400 2.5950 1.3700 ;
        RECT  2.3350 0.9400 2.5950 1.0900 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.4900 2.9550 1.6100 ;
        RECT  2.8350 1.1050 2.9550 1.6100 ;
        RECT  0.6800 1.2800 1.0750 1.6100 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1550 1.4650 3.4100 1.7250 ;
        RECT  0.4100 1.7300 3.3800 1.8500 ;
        RECT  3.1550 1.4650 3.3800 1.8500 ;
        RECT  3.1550 1.2200 3.2750 1.8500 ;
        RECT  0.4100 1.2200 0.5300 1.8500 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7350 0.4000 5.8550 0.9150 ;
        RECT  5.5550 0.7950 5.8550 0.9150 ;
        RECT  3.9950 0.9100 5.6750 1.0300 ;
        RECT  5.5350 1.3900 5.6550 2.2100 ;
        RECT  3.8550 1.3900 5.6550 1.5100 ;
        RECT  4.9350 1.1750 5.1500 1.5100 ;
        RECT  4.9350 0.9100 5.0550 1.5100 ;
        RECT  4.8950 0.4000 5.0150 1.0300 ;
        RECT  4.6950 1.3900 4.8150 2.2100 ;
        RECT  3.9950 0.4000 4.1150 1.0300 ;
        RECT  3.8550 1.3900 3.9750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.3150 -0.1800 5.4350 0.7900 ;
        RECT  4.4750 -0.1800 4.5950 0.7900 ;
        RECT  3.5150 0.4600 3.7550 0.5800 ;
        RECT  3.5150 -0.1800 3.6350 0.5800 ;
        RECT  2.6750 0.4600 2.9150 0.5800 ;
        RECT  2.6750 -0.1800 2.7950 0.5800 ;
        RECT  1.8350 0.4600 2.0750 0.5800 ;
        RECT  1.8350 -0.1800 1.9550 0.5800 ;
        RECT  0.9950 0.4600 1.2350 0.5800 ;
        RECT  0.9950 -0.1800 1.1150 0.5800 ;
        RECT  0.2150 -0.1800 0.3350 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1150 1.6300 5.2350 2.7900 ;
        RECT  4.2750 1.6300 4.3950 2.7900 ;
        RECT  3.3150 2.2100 3.5550 2.7900 ;
        RECT  0.4150 1.9700 0.5350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8150 1.2700 3.6500 1.2700 3.6500 2.0900 2.1750 2.0900 2.1750 2.1500 1.9350 2.1500
                 1.9350 1.9700 3.5300 1.9700 3.5300 0.8200 0.6950 0.8200 0.6950 0.7700 0.5750 0.7700
                 0.5750 0.6500 0.8150 0.6500 0.8150 0.7000 1.4150 0.7000 1.4150 0.6500 1.6550 0.6500
                 1.6550 0.7000 2.2550 0.7000 2.2550 0.6500 2.4950 0.6500 2.4950 0.7000 3.0950 0.7000
                 3.0950 0.6500 3.3350 0.6500 3.3350 0.7000 3.6500 0.7000 3.6500 1.1500 4.8150 1.1500 ;
    END
END OR4X6

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5150 1.0250 1.9600 1.1450 ;
        RECT  1.8100 0.8850 1.9600 1.1450 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0300 0.5100 1.4850 ;
        RECT  0.3600 1.0000 0.4800 1.4850 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0500 0.8200 1.4850 ;
        RECT  0.7000 1.0250 0.8200 1.4850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0350 1.1050 1.1550 1.4600 ;
        RECT  0.9400 1.1350 1.0900 1.4850 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0750 0.5900 3.1950 0.8300 ;
        RECT  2.0550 1.5050 3.1750 1.6250 ;
        RECT  3.0750 0.5900 3.1750 1.6250 ;
        RECT  2.8950 1.5050 3.1200 1.7250 ;
        RECT  2.9700 1.4650 3.1750 1.6250 ;
        RECT  3.0550 0.7100 3.1200 1.7250 ;
        RECT  2.2350 0.7600 3.1750 0.8800 ;
        RECT  2.8950 1.5050 3.0150 2.2100 ;
        RECT  2.2350 0.5900 2.3550 0.8800 ;
        RECT  2.0550 1.5050 2.1750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.4950 -0.1800 3.6150 0.6400 ;
        RECT  2.6550 -0.1800 2.7750 0.6400 ;
        RECT  1.8150 -0.1800 1.9350 0.6400 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.3150 1.5600 3.4350 2.7900 ;
        RECT  2.4750 1.7450 2.5950 2.7900 ;
        RECT  1.6350 1.5600 1.7550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.9350 1.3450 2.8500 1.3450 2.8500 1.3850 1.3950 1.3850 1.3950 1.7250 0.3400 1.7250
                 0.3400 2.2100 0.2200 2.2100 0.2200 1.6050 1.2750 1.6050 1.2750 0.8800 0.5550 0.8800
                 0.5550 0.5900 0.6750 0.5900 0.6750 0.7600 1.3950 0.7600 1.3950 0.5900 1.5150 0.5900
                 1.5150 0.8800 1.3950 0.8800 1.3950 1.2650 2.7300 1.2650 2.7300 1.1050 2.9350 1.1050 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9200 2.0150 1.1200 ;
        RECT  1.7550 0.8900 1.8750 1.2400 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3100 1.1750 0.5300 1.4350 ;
        RECT  0.3350 1.0600 0.5300 1.4350 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0350 0.8200 1.4400 ;
        RECT  0.7000 1.0200 0.8200 1.4400 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2550 1.0800 1.3750 1.3200 ;
        RECT  0.9400 1.1750 1.3750 1.2950 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.1750 2.5400 1.4350 ;
        RECT  2.4150 0.6800 2.5350 1.4350 ;
        RECT  2.3350 1.2950 2.4550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.8350 -0.1800 2.9550 0.7300 ;
        RECT  1.9950 -0.1800 2.1150 0.7300 ;
        RECT  1.0350 -0.1800 1.1550 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.9000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.7550 1.5600 2.8750 2.7900 ;
        RECT  1.9150 1.6000 2.0350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2150 1.4800 1.6350 1.4800 1.6350 1.6800 0.3400 1.6800 0.3400 1.8000 0.2200 1.8000
                 0.2200 1.5600 1.5150 1.5600 1.5150 0.9000 0.5550 0.9000 0.5550 0.6600 0.6750 0.6600
                 0.6750 0.7800 1.5150 0.7800 1.5150 0.6600 1.6350 0.6600 1.6350 1.3600 2.0950 1.3600
                 2.0950 1.2400 2.2150 1.2400 ;
    END
END OR4X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.8350 1.9600 1.1500 ;
        RECT  1.6550 1.0300 1.9300 1.1800 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2850 1.1750 0.5250 1.4350 ;
        RECT  0.1850 1.2600 0.4050 1.5000 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 1.0200 0.8450 1.2850 ;
        RECT  0.6450 1.1650 0.8200 1.4450 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2400 1.2950 1.5250 ;
        RECT  0.9700 1.4050 1.2950 1.5250 ;
        RECT  0.9400 1.4650 1.0900 1.7250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3550 1.1750 2.5400 1.4350 ;
        RECT  2.3550 0.6600 2.4750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.9350 -0.1800 2.0550 0.7100 ;
        RECT  1.0350 -0.1800 1.1550 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.9000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.9350 1.5600 2.0550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2350 1.4200 1.5350 1.4200 1.5350 1.9650 0.4750 1.9650 0.4750 1.7000 0.5950 1.7000
                 0.5950 1.8450 1.4150 1.8450 1.4150 0.9000 0.5550 0.9000 0.5550 0.6600 0.6750 0.6600
                 0.6750 0.7800 1.4550 0.7800 1.4550 0.6600 1.5750 0.6600 1.5750 0.9000 1.5350 0.9000
                 1.5350 1.3000 2.2350 1.3000 ;
    END
END OR4X1

MACRO OR3XL
    CLASS CORE ;
    FOREIGN OR3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0000 0.5100 1.4550 ;
        RECT  0.3600 1.0000 0.4800 1.4800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6950 1.0200 0.8150 1.4550 ;
        RECT  0.6500 1.0200 0.8150 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2050 1.4350 1.4200 ;
        RECT  1.1750 1.0400 1.2950 1.4200 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6550 1.2950 1.9600 1.4350 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        RECT  1.8150 0.4000 1.9350 0.6400 ;
        RECT  1.8100 0.5200 1.9300 1.4350 ;
        RECT  1.6550 1.2950 1.7750 1.6600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.2350 1.5400 1.3550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6150 1.0400 1.4950 1.0400 1.4950 0.9200 1.0550 0.9200 1.0550 1.7200 0.1550 1.7200
                 0.1550 1.6000 0.9350 1.6000 0.9350 0.8800 0.1350 0.8800 0.1350 0.4000 0.2550 0.4000
                 0.2550 0.7600 0.9750 0.7600 0.9750 0.4000 1.0950 0.4000 1.0950 0.8000 1.6150 0.8000 ;
    END
END OR3XL

MACRO OR3X8
    CLASS CORE ;
    FOREIGN OR3X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6100 0.8200 2.7300 1.1700 ;
        RECT  0.3900 0.8200 2.7300 0.9400 ;
        RECT  0.3900 0.8200 0.5100 1.1500 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0600 2.3900 1.3000 ;
        RECT  2.1000 1.0600 2.2500 1.4350 ;
        RECT  1.0300 1.0600 2.3900 1.1800 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.3000 1.7900 1.4200 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.5500 1.3000 1.6700 1.7250 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9500 0.7150 6.1900 0.8350 ;
        RECT  3.5500 0.7650 6.0700 0.8850 ;
        RECT  5.8100 1.4700 5.9300 2.2100 ;
        RECT  5.6300 1.4700 5.9300 1.5900 ;
        RECT  5.6300 1.2750 5.7500 1.5900 ;
        RECT  3.2900 1.2750 5.7500 1.3950 ;
        RECT  5.1900 0.7650 5.4400 1.1450 ;
        RECT  5.1900 0.7650 5.3100 1.3950 ;
        RECT  5.1700 0.6450 5.2900 0.8850 ;
        RECT  4.9700 1.2750 5.2700 1.5900 ;
        RECT  4.9700 1.2750 5.0900 2.2100 ;
        RECT  4.2700 0.7150 4.5100 0.8850 ;
        RECT  4.1300 1.2750 4.2500 2.2100 ;
        RECT  3.4300 0.7150 3.6700 0.8350 ;
        RECT  3.2900 1.2750 3.4100 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.5900 -0.1800 5.7100 0.6450 ;
        RECT  4.7500 -0.1800 4.8700 0.6450 ;
        RECT  3.9100 -0.1800 4.0300 0.6450 ;
        RECT  2.9500 0.3400 3.1900 0.4600 ;
        RECT  2.9500 -0.1800 3.0700 0.4600 ;
        RECT  1.9900 0.3400 2.2300 0.4600 ;
        RECT  1.9900 -0.1800 2.1100 0.4600 ;
        RECT  1.0300 0.3400 1.2700 0.4600 ;
        RECT  1.0300 -0.1800 1.1500 0.4600 ;
        RECT  0.1900 -0.1800 0.3100 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.3900 1.5150 5.5100 2.7900 ;
        RECT  4.5500 1.5150 4.6700 2.7900 ;
        RECT  3.7100 1.5150 3.8300 2.7900 ;
        RECT  2.8700 1.7950 2.9900 2.7900 ;
        RECT  0.6100 1.5600 0.7300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.0700 1.1550 2.9700 1.1550 2.9700 1.6750 1.9100 1.6750 1.9100 2.2100 1.7900 2.2100
                 1.7900 1.5550 2.8500 1.5550 2.8500 0.7000 0.5500 0.7000 0.5500 0.5800 2.9700 0.5800
                 2.9700 1.0350 5.0700 1.0350 ;
    END
END OR3X8

MACRO OR3X6
    CLASS CORE ;
    FOREIGN OR3X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6700 0.8200 2.7900 1.1700 ;
        RECT  0.3900 0.8200 2.7900 0.9400 ;
        RECT  0.3900 0.8200 0.5100 1.1500 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0600 2.3900 1.3000 ;
        RECT  2.1000 1.0600 2.2500 1.4350 ;
        RECT  1.0300 1.0600 2.3900 1.1800 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.3000 1.7900 1.4200 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.5500 1.3000 1.6700 1.7250 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4900 0.9300 5.3500 1.0500 ;
        RECT  5.2300 0.4000 5.3500 1.0500 ;
        RECT  5.0300 1.4100 5.1500 2.2100 ;
        RECT  3.3500 1.4100 5.1500 1.5300 ;
        RECT  4.4100 0.8850 4.5700 1.1450 ;
        RECT  4.4100 0.7950 4.5300 1.5300 ;
        RECT  4.3900 0.4000 4.5100 1.0500 ;
        RECT  4.1900 1.4100 4.3100 2.2100 ;
        RECT  3.4900 0.4000 3.6100 1.0500 ;
        RECT  3.3500 1.4100 3.4700 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.8100 -0.1800 4.9300 0.8100 ;
        RECT  3.9700 -0.1800 4.0900 0.8100 ;
        RECT  2.9500 0.3400 3.1900 0.4600 ;
        RECT  2.9500 -0.1800 3.0700 0.4600 ;
        RECT  1.9900 0.3400 2.2300 0.4600 ;
        RECT  1.9900 -0.1800 2.1100 0.4600 ;
        RECT  1.0300 0.3400 1.2700 0.4600 ;
        RECT  1.0300 -0.1800 1.1500 0.4600 ;
        RECT  0.1900 -0.1800 0.3100 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.6100 1.6500 4.7300 2.7900 ;
        RECT  3.7700 1.6500 3.8900 2.7900 ;
        RECT  2.9300 1.7950 3.0500 2.7900 ;
        RECT  0.6100 1.5600 0.7300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.2900 1.2900 3.0300 1.2900 3.0300 1.6750 1.9100 1.6750 1.9100 2.2100 1.7900 2.2100
                 1.7900 1.5550 2.9100 1.5550 2.9100 0.7000 0.5500 0.7000 0.5500 0.5800 3.0300 0.5800
                 3.0300 1.1700 4.2900 1.1700 ;
    END
END OR3X6

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0000 0.5100 1.4500 ;
        RECT  0.3600 1.0000 0.4800 1.4750 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7500 1.0000 0.8700 1.3450 ;
        RECT  0.6500 1.0900 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.3700 1.3800 1.7250 ;
        RECT  1.2300 1.2300 1.3500 1.7250 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.8850 3.1200 1.1450 ;
        RECT  2.7100 0.8850 3.1200 1.0050 ;
        RECT  2.5700 1.5600 2.8300 1.6800 ;
        RECT  2.7100 0.7100 2.8300 1.6800 ;
        RECT  2.6700 0.5900 2.7900 0.8300 ;
        RECT  1.7300 1.3200 2.8300 1.4400 ;
        RECT  2.5700 1.5600 2.6900 2.2100 ;
        RECT  1.8900 0.7100 2.8300 0.8300 ;
        RECT  1.7700 0.6500 2.0100 0.7700 ;
        RECT  1.7300 1.3200 1.8500 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  3.0900 -0.1800 3.2100 0.6400 ;
        RECT  2.1900 0.4600 2.4300 0.5800 ;
        RECT  2.1900 -0.1800 2.3100 0.5800 ;
        RECT  1.4100 -0.1800 1.5300 0.6400 ;
        RECT  0.5700 -0.1800 0.6900 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.9900 1.5600 3.1100 2.7900 ;
        RECT  2.1500 1.5600 2.2700 2.7900 ;
        RECT  1.3100 1.8450 1.4300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.5900 1.1100 1.1100 1.1100 1.1100 1.7150 0.3900 1.7150 0.3900 2.2100 0.2700 2.2100
                 0.2700 1.5950 0.9900 1.5950 0.9900 0.8800 0.1500 0.8800 0.1500 0.5900 0.2700 0.5900
                 0.2700 0.7600 0.9900 0.7600 0.9900 0.5900 1.1100 0.5900 1.1100 0.9900 2.5900 0.9900 ;
    END
END OR3X4

MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0000 0.5100 1.4550 ;
        RECT  0.3750 1.0000 0.4950 1.4850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6950 1.0050 0.8150 1.4650 ;
        RECT  0.6500 1.0000 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 0.9400 1.4350 1.2000 ;
        RECT  1.1750 0.9400 1.4150 1.2200 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8150 1.0250 2.2500 1.1450 ;
        RECT  2.1000 0.8850 2.2500 1.1450 ;
        RECT  1.8150 0.5900 1.9350 1.3900 ;
        RECT  1.7150 1.2700 1.8350 1.9900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  2.2350 -0.1800 2.3550 0.6400 ;
        RECT  1.3350 0.4600 1.5750 0.5800 ;
        RECT  1.3350 -0.1800 1.4550 0.5800 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  2.1350 1.3400 2.2550 2.7900 ;
        RECT  1.2950 1.3400 1.4150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6950 1.1500 1.5750 1.1500 1.5750 0.8200 1.0550 0.8200 1.0550 1.7250 0.1550 1.7250
                 0.1550 1.6050 0.9350 1.6050 0.9350 0.8800 0.1350 0.8800 0.1350 0.4000 0.2550 0.4000
                 0.2550 0.7600 0.9350 0.7600 0.9350 0.7000 0.9750 0.7000 0.9750 0.4000 1.0950 0.4000
                 1.0950 0.7000 1.6950 0.7000 ;
    END
END OR3X2

MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0000 0.5100 1.4550 ;
        RECT  0.3750 1.0000 0.4950 1.4850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6950 1.0000 0.8150 1.4600 ;
        RECT  0.6500 1.0000 0.8150 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 0.9400 1.4350 1.2100 ;
        RECT  1.1750 0.9400 1.4150 1.2200 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.8850 1.9600 1.1450 ;
        RECT  1.8150 0.5900 1.9350 1.1450 ;
        RECT  1.7950 1.1450 1.9300 1.2650 ;
        RECT  1.7950 1.1450 1.9150 1.9900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3350 0.4600 1.5750 0.5800 ;
        RECT  1.3350 -0.1800 1.4550 0.5800 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.3750 1.3400 1.4950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6750 1.1700 1.5550 1.1700 1.5550 0.8200 1.0550 0.8200 1.0550 1.7250 0.1550 1.7250
                 0.1550 1.6050 0.9350 1.6050 0.9350 0.8800 0.1350 0.8800 0.1350 0.4000 0.2550 0.4000
                 0.2550 0.7600 0.9350 0.7600 0.9350 0.7000 0.9750 0.7000 0.9750 0.4000 1.0950 0.4000
                 1.0950 0.7000 1.6750 0.7000 ;
    END
END OR3X1

MACRO OR2XL
    CLASS CORE ;
    FOREIGN OR2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.3950 1.3200 ;
        RECT  0.2750 1.0800 0.3950 1.3200 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.3900 1.0900 1.7250 ;
        RECT  0.8150 1.3900 1.0900 1.6250 ;
        RECT  0.8150 1.2900 0.9350 1.6250 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4850 0.6800 1.6050 0.9200 ;
        RECT  1.3950 0.8000 1.5150 1.9650 ;
        RECT  1.2300 1.4650 1.5150 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  1.0350 -0.1800 1.1550 0.4000 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.8450 1.0950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.2550 1.2700 1.1350 1.2700 1.1350 1.1700 0.6750 1.1700 0.6750 1.9050 0.2750 1.9050
                 0.2750 1.7850 0.5550 1.7850 0.5550 0.6800 0.6750 0.6800 0.6750 1.0500 1.1350 1.0500
                 1.1350 1.0300 1.2550 1.0300 ;
    END
END OR2XL

MACRO OR2X8
    CLASS CORE ;
    FOREIGN OR2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0550 1.6350 1.1750 ;
        RECT  0.3600 1.1750 0.5600 1.2950 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.2950 1.0150 1.4150 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.2950 0.8000 1.7250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6950 0.7150 4.9350 0.8350 ;
        RECT  2.2950 0.7650 4.8150 0.8850 ;
        RECT  4.6150 1.4700 4.7350 2.2100 ;
        RECT  4.4350 1.4700 4.7350 1.5900 ;
        RECT  4.4350 1.2750 4.5550 1.5900 ;
        RECT  2.0950 1.2750 4.5550 1.3950 ;
        RECT  3.9350 0.7650 4.2800 1.1450 ;
        RECT  3.9350 0.7650 4.0550 1.3950 ;
        RECT  3.9150 0.6450 4.0350 0.8850 ;
        RECT  3.7750 1.2750 3.8950 2.2100 ;
        RECT  3.0150 0.7150 3.2550 0.8850 ;
        RECT  2.9350 1.2750 3.0550 2.2100 ;
        RECT  2.1750 0.7150 2.4150 0.8350 ;
        RECT  2.0950 1.2750 2.2150 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  4.3350 -0.1800 4.4550 0.6450 ;
        RECT  3.4950 -0.1800 3.6150 0.6450 ;
        RECT  2.6550 -0.1800 2.7750 0.6450 ;
        RECT  1.8150 -0.1800 1.9350 0.6950 ;
        RECT  0.9750 -0.1800 1.0950 0.6950 ;
        RECT  0.1350 -0.1800 0.2550 0.6950 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  4.1950 1.5150 4.3150 2.7900 ;
        RECT  3.3550 1.5150 3.4750 2.7900 ;
        RECT  2.5150 1.5150 2.6350 2.7900 ;
        RECT  1.6750 1.5550 1.7950 2.7900 ;
        RECT  0.3350 1.5550 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.8150 1.1550 1.8750 1.1550 1.8750 1.4150 1.2550 1.4150 1.2550 1.6750 1.0950 1.6750
                 1.0950 2.2050 0.9750 2.2050 0.9750 1.5550 1.1350 1.5550 1.1350 1.2950 1.7550 1.2950
                 1.7550 0.9350 0.5550 0.9350 0.5550 0.6450 0.6750 0.6450 0.6750 0.8150 1.3950 0.8150
                 1.3950 0.6450 1.5150 0.6450 1.5150 0.8150 1.8750 0.8150 1.8750 1.0350 3.8150 1.0350 ;
    END
END OR2X8

MACRO OR2X6
    CLASS CORE ;
    FOREIGN OR2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0600 1.6350 1.1800 ;
        RECT  0.3600 1.1750 0.5600 1.3000 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.3000 1.0150 1.4200 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.3000 0.8000 1.7250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2350 0.9100 4.0950 1.0300 ;
        RECT  3.9750 0.4000 4.0950 1.0300 ;
        RECT  3.7750 1.3900 3.8950 2.2100 ;
        RECT  2.0950 1.3900 3.8950 1.5100 ;
        RECT  3.1750 0.8850 3.4100 1.1450 ;
        RECT  3.1750 0.7950 3.2950 1.5100 ;
        RECT  3.1350 0.4000 3.2550 1.0300 ;
        RECT  2.9350 1.3900 3.0550 2.2100 ;
        RECT  2.2350 0.4000 2.3550 1.0300 ;
        RECT  2.0950 1.3900 2.2150 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.5550 -0.1800 3.6750 0.7900 ;
        RECT  2.7150 -0.1800 2.8350 0.7900 ;
        RECT  1.8150 -0.1800 1.9350 0.7000 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.3550 1.6300 3.4750 2.7900 ;
        RECT  2.5150 1.6300 2.6350 2.7900 ;
        RECT  1.6750 1.5600 1.7950 2.7900 ;
        RECT  0.3350 1.5600 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0550 1.2700 1.8750 1.2700 1.8750 1.4400 1.2550 1.4400 1.2550 1.6800 1.0950 1.6800
                 1.0950 2.2100 0.9750 2.2100 0.9750 1.5600 1.1350 1.5600 1.1350 1.3200 1.7550 1.3200
                 1.7550 0.9400 0.5550 0.9400 0.5550 0.5900 0.6750 0.5900 0.6750 0.8200 1.3950 0.8200
                 1.3950 0.5900 1.5150 0.5900 1.5150 0.8200 1.8750 0.8200 1.8750 1.1500 3.0550 1.1500 ;
    END
END OR2X6

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.9500 0.5100 1.1900 ;
        RECT  0.0700 0.9500 0.5100 1.0700 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.4500 1.0900 1.7250 ;
        RECT  0.9300 1.3550 1.0600 1.4750 ;
        RECT  0.9300 1.2200 1.0500 1.4750 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.3900 0.7400 2.5100 1.6800 ;
        RECT  2.3500 1.5600 2.4700 2.2100 ;
        RECT  1.5100 1.3200 2.5100 1.4400 ;
        RECT  1.5700 0.7400 2.5100 0.8600 ;
        RECT  2.3500 0.6200 2.4700 0.8600 ;
        RECT  1.4500 0.6900 1.6900 0.8100 ;
        RECT  1.5100 1.3200 1.6300 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.7700 -0.1800 2.8900 0.6800 ;
        RECT  1.8700 0.5000 2.1100 0.6200 ;
        RECT  1.8700 -0.1800 1.9900 0.6200 ;
        RECT  1.0900 -0.1800 1.2100 0.6800 ;
        RECT  0.2500 -0.1800 0.3700 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.7700 1.5600 2.8900 2.7900 ;
        RECT  1.9300 1.5600 2.0500 2.7900 ;
        RECT  1.0900 1.8450 1.2100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2700 1.1500 2.0300 1.1500 2.0300 1.1000 1.8500 1.1000 1.8500 1.1500 1.6100 1.1500
                 1.6100 1.1000 0.7900 1.1000 0.7900 1.4300 0.5700 1.4300 0.5700 2.2100 0.4500 2.2100
                 0.4500 1.3100 0.6700 1.3100 0.6700 0.6300 0.7900 0.6300 0.7900 0.9800 2.1500 0.9800
                 2.1500 1.0300 2.2700 1.0300 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2350 0.9800 0.3550 1.2200 ;
        RECT  0.0700 0.9800 0.3550 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.2150 1.1450 1.3800 ;
        RECT  0.7750 1.2000 0.8950 1.4750 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5050 0.8850 1.6700 1.1450 ;
        RECT  1.3550 1.3600 1.6250 1.4800 ;
        RECT  1.5050 0.7200 1.6250 1.4800 ;
        RECT  1.3550 0.7200 1.6250 0.8400 ;
        RECT  1.3550 1.3600 1.4750 2.2100 ;
        RECT  1.3550 0.6000 1.4750 0.8400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  1.7750 -0.1800 1.8950 0.7300 ;
        RECT  0.8750 0.7200 1.1150 0.8400 ;
        RECT  0.8750 -0.1800 0.9950 0.8400 ;
        RECT  0.1350 -0.1800 0.2550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.7750 1.5600 1.8950 2.7900 ;
        RECT  0.9350 1.5950 1.0550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.3850 1.2400 1.2650 1.2400 1.2650 1.0800 0.6350 1.0800 0.6350 1.4600 0.4150 1.4600
                 0.4150 1.7400 0.1750 1.7400 0.1750 1.6200 0.2950 1.6200 0.2950 1.3400 0.5150 1.3400
                 0.5150 0.6600 0.6350 0.6600 0.6350 0.9600 1.3850 0.9600 ;
    END
END OR2X2

MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.0250 0.4250 1.2650 ;
        RECT  0.0700 1.0250 0.4250 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8450 1.1750 1.1450 1.3800 ;
        RECT  0.8450 1.0700 0.9650 1.4300 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5050 0.8850 1.6700 1.1450 ;
        RECT  1.5050 0.5900 1.6250 1.4800 ;
        RECT  1.4850 1.3600 1.6050 2.2000 ;
        RECT  1.4850 0.4700 1.6050 0.7100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  1.0050 0.5300 1.2450 0.6500 ;
        RECT  1.0050 -0.1800 1.1250 0.6500 ;
        RECT  0.1350 -0.1800 0.2550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.0650 1.5500 1.1850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.3850 1.2400 1.2650 1.2400 1.2650 0.9500 0.7050 0.9500 0.7050 1.5050 0.5450 1.5050
                 0.5450 1.7300 0.3050 1.7300 0.3050 1.6100 0.4250 1.6100 0.4250 1.3850 0.5850 1.3850
                 0.5850 0.6600 0.7050 0.6600 0.7050 0.8300 1.3850 0.8300 ;
    END
END OR2X1

MACRO OAI33XL
    CLASS CORE ;
    FOREIGN OAI33XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3700 1.1400 2.6100 1.3450 ;
        RECT  2.3900 1.0800 2.5400 1.4750 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1050 2.2500 1.5600 ;
        RECT  2.1000 1.0800 2.2200 1.5600 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.1750 1.3800 1.6750 ;
        RECT  1.2300 1.1750 1.3800 1.6450 ;
        END
    END A2
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4200 1.2400 0.5400 1.6200 ;
        RECT  0.0700 1.3150 0.5400 1.4350 ;
        RECT  0.0700 1.0600 0.2200 1.4350 ;
        END
    END A0
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.3350 1.8600 1.4850 ;
        RECT  1.5200 1.1400 1.6700 1.4550 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1400 1.0900 1.6100 ;
        RECT  0.9400 1.1400 1.0600 1.6400 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2592  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7800 0.5400 2.9000 0.7800 ;
        RECT  1.5200 1.6800 2.8500 1.8000 ;
        RECT  2.6800 1.4650 2.8500 1.8000 ;
        RECT  2.7300 0.6600 2.8500 1.8000 ;
        RECT  2.0000 0.8400 2.8500 0.9600 ;
        RECT  2.0000 0.6000 2.1200 0.9600 ;
        RECT  1.8800 0.6000 2.1200 0.7200 ;
        RECT  1.5200 1.6800 1.6400 2.0400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  1.1000 -0.1800 1.2200 0.7800 ;
        RECT  0.2600 -0.1800 0.3800 0.7800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.5800 1.9200 2.7000 2.7900 ;
        RECT  0.4600 1.9200 0.5800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.5400 0.7200 2.3000 0.7200 2.3000 0.4800 1.6400 0.4800 1.6400 1.0200 0.6800 1.0200
                 0.6800 0.5400 0.8000 0.5400 0.8000 0.9000 1.5200 0.9000 1.5200 0.3600 2.4200 0.3600
                 2.4200 0.6000 2.5400 0.6000 ;
    END
END OAI33XL

MACRO OAI33X4
    CLASS CORE ;
    FOREIGN OAI33X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8450 1.2600 8.8550 1.3800 ;
        RECT  7.8450 1.2300 8.1050 1.3800 ;
        RECT  7.9550 1.0000 8.0750 1.3800 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1750 1.6700 1.4350 ;
        RECT  1.5350 0.9400 1.6550 1.4350 ;
        RECT  0.8950 1.2800 1.6700 1.4000 ;
        RECT  0.7750 1.3000 1.0150 1.4200 ;
        END
    END A0
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.5350 1.2200 5.0950 1.3400 ;
        RECT  4.6550 1.2200 4.9150 1.3800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.1750 3.4100 1.4350 ;
        RECT  3.2600 0.9400 3.3800 1.4350 ;
        RECT  2.4350 1.2800 3.4100 1.4000 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.2150 1.2200 6.7750 1.3400 ;
        RECT  6.3950 1.2200 6.6550 1.3800 ;
        END
    END B2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6550 1.2600 10.5550 1.3800 ;
        RECT  9.6550 1.2300 10.1350 1.3800 ;
        RECT  9.6550 1.0000 9.7750 1.3800 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.8136  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1550 0.6500 10.3950 0.7700 ;
        RECT  5.9550 0.7600 10.2750 0.8800 ;
        RECT  9.3150 0.6500 9.5550 0.8800 ;
        RECT  8.4750 0.6500 8.7150 0.8800 ;
        RECT  7.6350 0.6500 7.8750 0.8800 ;
        RECT  7.2750 1.5000 7.3950 2.0100 ;
        RECT  3.9150 1.5000 7.3950 1.6200 ;
        RECT  6.7950 0.6500 7.0350 0.8800 ;
        RECT  6.4350 1.5000 6.5550 2.0100 ;
        RECT  5.9550 0.6500 6.1950 0.8800 ;
        RECT  4.2150 0.9800 6.0750 1.1000 ;
        RECT  5.9550 0.6500 6.0750 1.1000 ;
        RECT  5.5950 1.5000 5.7150 2.1500 ;
        RECT  4.7550 1.5000 4.8750 2.0100 ;
        RECT  4.2150 0.9800 4.3350 1.6200 ;
        RECT  4.0750 1.2300 4.3350 1.3800 ;
        RECT  3.9150 1.5000 4.0350 2.0100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  5.1150 0.4600 5.3550 0.5800 ;
        RECT  5.1150 -0.1800 5.2350 0.5800 ;
        RECT  4.2750 0.4600 4.5150 0.5800 ;
        RECT  4.2750 -0.1800 4.3950 0.5800 ;
        RECT  3.4350 0.4600 3.6750 0.5800 ;
        RECT  3.4350 -0.1800 3.5550 0.5800 ;
        RECT  2.5950 0.4600 2.8350 0.5800 ;
        RECT  2.5950 -0.1800 2.7150 0.5800 ;
        RECT  1.7550 0.4600 1.9950 0.5800 ;
        RECT  1.7550 -0.1800 1.8750 0.5800 ;
        RECT  0.9150 0.4600 1.1550 0.5800 ;
        RECT  0.9150 -0.1800 1.0350 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.6350 1.7400 10.7550 2.7900 ;
        RECT  9.7950 1.7400 9.9150 2.7900 ;
        RECT  1.3950 1.7950 1.5150 2.7900 ;
        RECT  0.5550 1.7950 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.1750 2.2100 11.0550 2.2100 11.0550 1.6200 10.3350 1.6200 10.3350 2.2100
                 10.2150 2.2100 10.2150 1.6200 9.4950 1.6200 9.4950 2.2100 9.3750 2.2100 9.3750 1.6200
                 8.6550 1.6200 8.6550 2.0100 8.5350 2.0100 8.5350 1.6200 7.8150 1.6200 7.8150 2.0100
                 7.6950 2.0100 7.6950 1.5000 11.1750 1.5000 ;
        POLYGON  10.7550 0.6500 10.6350 0.6500 10.6350 0.5300 9.9150 0.5300 9.9150 0.6400 9.7950 0.6400
                 9.7950 0.5300 9.0750 0.5300 9.0750 0.6400 8.9550 0.6400 8.9550 0.5300 8.2350 0.5300
                 8.2350 0.6400 8.1150 0.6400 8.1150 0.5300 7.3950 0.5300 7.3950 0.6400 7.2750 0.6400
                 7.2750 0.5300 6.5550 0.5300 6.5550 0.6400 6.4350 0.6400 6.4350 0.5300 5.7150 0.5300
                 5.7150 0.8200 0.5550 0.8200 0.5550 0.5800 0.6750 0.5800 0.6750 0.7000 1.3950 0.7000
                 1.3950 0.5800 1.5150 0.5800 1.5150 0.7000 2.2350 0.7000 2.2350 0.5800 2.3550 0.5800
                 2.3550 0.7000 3.0750 0.7000 3.0750 0.5800 3.1950 0.5800 3.1950 0.7000 3.9150 0.7000
                 3.9150 0.5800 4.0350 0.5800 4.0350 0.7000 4.7550 0.7000 4.7550 0.5800 4.8750 0.5800
                 4.8750 0.7000 5.5950 0.7000 5.5950 0.4100 6.4350 0.4100 6.4350 0.4000 6.5550 0.4000
                 6.5550 0.4100 7.2750 0.4100 7.2750 0.4000 7.3950 0.4000 7.3950 0.4100 8.1150 0.4100
                 8.1150 0.4000 8.2350 0.4000 8.2350 0.4100 8.9550 0.4100 8.9550 0.4000 9.0750 0.4000
                 9.0750 0.4100 9.7950 0.4100 9.7950 0.4000 9.9150 0.4000 9.9150 0.4100 10.7550 0.4100 ;
        POLYGON  9.0750 2.2500 6.0150 2.2500 6.0150 1.7400 6.1350 1.7400 6.1350 2.1300 6.8550 2.1300
                 6.8550 1.7400 6.9750 1.7400 6.9750 2.1300 8.1150 2.1300 8.1150 1.7400 8.2350 1.7400
                 8.2350 2.1300 8.9550 2.1300 8.9550 1.7400 9.0750 1.7400 ;
        POLYGON  5.2950 2.2500 2.2350 2.2500 2.2350 1.7950 2.3550 1.7950 2.3550 2.1300 3.0750 2.1300
                 3.0750 1.7950 3.1950 1.7950 3.1950 2.1300 4.3350 2.1300 4.3350 1.7400 4.4550 1.7400
                 4.4550 2.1300 5.1750 2.1300 5.1750 1.7400 5.2950 1.7400 ;
        POLYGON  3.6150 2.0100 3.4950 2.0100 3.4950 1.6750 2.7750 1.6750 2.7750 2.0100 2.6550 2.0100
                 2.6550 1.6750 1.9350 1.6750 1.9350 2.2100 1.8150 2.2100 1.8150 1.6750 1.0950 1.6750
                 1.0950 2.2100 0.9750 2.2100 0.9750 1.6750 0.2550 1.6750 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.5550 3.6150 1.5550 ;
    END
END OAI33X4

MACRO OAI33X2
    CLASS CORE ;
    FOREIGN OAI33X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0086  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0750 0.6600 8.3750 0.7800 ;
        RECT  8.2550 0.5400 8.3750 0.7800 ;
        RECT  7.3550 0.8550 8.1950 0.9750 ;
        RECT  8.0750 0.6600 8.1950 0.9750 ;
        RECT  1.4550 1.8450 7.9950 1.9650 ;
        RECT  7.8750 0.8550 7.9950 1.9650 ;
        RECT  7.3550 0.6000 7.5950 0.7200 ;
        RECT  4.8200 0.7900 7.4750 0.9100 ;
        RECT  7.3550 0.6000 7.4750 0.9750 ;
        RECT  6.4550 0.6000 6.6950 0.9100 ;
        RECT  5.6150 0.6000 5.8550 0.9100 ;
        RECT  4.6550 0.6500 5.0150 0.8000 ;
        RECT  4.7750 0.6000 5.0150 0.8000 ;
        END
    END Y
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2175  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4350 0.9700 2.8150 1.0900 ;
        RECT  2.3350 0.9400 2.5950 1.0900 ;
        END
    END A0
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2175  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7400 1.0300 7.1750 1.1500 ;
        RECT  4.7400 1.0300 4.9550 1.2950 ;
        RECT  4.7100 1.1750 4.8600 1.4350 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2175  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 1.2300 3.7750 1.3500 ;
        RECT  3.4950 1.2300 3.7550 1.3800 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2175  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.1350 1.2700 7.4950 1.3900 ;
        RECT  5.1350 1.2700 5.2550 1.5350 ;
        RECT  5.0000 1.4650 5.2150 1.6550 ;
        RECT  5.0000 1.4650 5.1500 1.7250 ;
        RECT  5.0300 1.4150 5.2550 1.5350 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2175  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0750 1.5200 4.3350 1.6700 ;
        RECT  1.2950 1.5000 4.3150 1.6100 ;
        RECT  4.0750 1.4900 4.3150 1.6700 ;
        RECT  1.9450 1.5200 4.3350 1.6200 ;
        RECT  1.2950 1.4900 2.0650 1.6100 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2175  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6350 1.4400 7.7550 1.6800 ;
        RECT  5.4750 1.5100 7.7550 1.6300 ;
        RECT  5.5250 1.5100 5.7850 1.6700 ;
        END
    END B0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  3.8550 0.4600 4.0950 0.5800 ;
        RECT  3.8550 -0.1800 3.9750 0.5800 ;
        RECT  2.8950 0.4600 3.1350 0.5800 ;
        RECT  2.8950 -0.1800 3.0150 0.5800 ;
        RECT  1.9350 0.4600 2.1750 0.5800 ;
        RECT  1.9350 -0.1800 2.0550 0.5800 ;
        RECT  0.9750 0.4600 1.2150 0.5800 ;
        RECT  0.9750 -0.1800 1.0950 0.5800 ;
        RECT  0.1350 -0.1800 0.2550 0.7250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.7950 2.0850 8.0350 2.2050 ;
        RECT  7.7950 2.0850 7.9150 2.7900 ;
        RECT  5.6550 2.0850 5.8950 2.2050 ;
        RECT  5.6550 2.0850 5.7750 2.7900 ;
        RECT  2.4750 2.0850 2.7150 2.2050 ;
        RECT  2.4750 2.0850 2.5950 2.7900 ;
        RECT  0.3350 1.9700 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.9550 0.7350 7.8350 0.7350 7.8350 0.4800 7.1150 0.4800 7.1150 0.6700 6.8750 0.6700
                 6.8750 0.4800 6.2750 0.4800 6.2750 0.6700 6.0350 0.6700 6.0350 0.4800 5.4350 0.4800
                 5.4350 0.6700 5.1950 0.6700 5.1950 0.4800 4.5350 0.4800 4.5350 0.8200 0.5550 0.8200
                 0.5550 0.5350 0.6750 0.5350 0.6750 0.7000 1.5150 0.7000 1.5150 0.5350 1.6350 0.5350
                 1.6350 0.7000 2.4750 0.7000 2.4750 0.5350 2.5950 0.5350 2.5950 0.7000 3.4350 0.7000
                 3.4350 0.5350 3.5550 0.5350 3.5550 0.7000 4.4150 0.7000 4.4150 0.3600 7.9550 0.3600 ;
    END
END OAI33X2

MACRO OAI33X1
    CLASS CORE ;
    FOREIGN OAI33X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0100 2.5400 1.4650 ;
        RECT  2.3900 1.0100 2.5100 1.4950 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8850 1.0550 2.0500 1.2950 ;
        RECT  1.8100 1.1750 2.0050 1.4350 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.0400 1.3800 1.4950 ;
        RECT  1.2500 1.0100 1.3700 1.4950 ;
        END
    END A2
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0100 0.5100 1.4650 ;
        RECT  0.3600 1.0100 0.4800 1.4950 ;
        END
    END A0
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5700 1.0200 1.6900 1.4350 ;
        RECT  1.5200 1.0950 1.6700 1.4950 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1500 1.0900 1.4350 ;
        RECT  0.8300 1.0200 0.9500 1.2950 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4660  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6600 1.4650 2.8300 1.7250 ;
        RECT  1.8300 0.7700 2.7900 0.8900 ;
        RECT  2.6700 0.6000 2.7900 0.8900 ;
        RECT  1.4100 1.6150 2.7800 1.7350 ;
        RECT  2.6600 0.7700 2.7800 1.7350 ;
        RECT  1.8300 0.6000 1.9500 0.8900 ;
        RECT  1.4100 1.6150 1.5300 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  0.9900 -0.1800 1.1100 0.6500 ;
        RECT  0.1500 -0.1800 0.2700 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3700 1.8550 2.4900 2.7900 ;
        RECT  0.3500 1.6150 0.4700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3700 0.6500 2.2500 0.6500 2.2500 0.5300 2.0700 0.5300 2.0700 0.4800 1.5300 0.4800
                 1.5300 0.8900 0.5700 0.8900 0.5700 0.6000 0.6900 0.6000 0.6900 0.7700 1.4100 0.7700
                 1.4100 0.3600 2.1900 0.3600 2.1900 0.4100 2.3700 0.4100 ;
    END
END OAI33X1

MACRO OAI32XL
    CLASS CORE ;
    FOREIGN OAI32XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.1750 2.5400 1.4350 ;
        RECT  2.1650 1.1750 2.5400 1.2950 ;
        RECT  2.1650 1.0550 2.2850 1.2950 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.3600 1.2950 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.4650 2.2500 1.7250 ;
        RECT  1.8450 1.5350 2.2500 1.6550 ;
        RECT  1.8450 1.4150 1.9650 1.6550 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 1.1750 0.8200 1.6100 ;
        RECT  0.6500 1.1750 0.8200 1.5900 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.3400 0.5100 1.7550 ;
        RECT  0.3600 1.0300 0.4800 1.7550 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2370  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5850 1.1750 2.0000 1.2950 ;
        RECT  1.8800 0.6350 2.0000 1.2950 ;
        RECT  1.4650 1.5200 1.7250 1.6700 ;
        RECT  1.5850 1.1750 1.7050 1.9950 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  0.9800 0.6950 1.2200 0.8150 ;
        RECT  0.9800 -0.1800 1.1000 0.8150 ;
        RECT  0.2000 -0.1800 0.3200 0.8750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  2.3250 1.8750 2.4450 2.7900 ;
        RECT  0.2000 1.8750 0.3200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4200 0.8750 2.3000 0.8750 2.3000 0.5150 1.5800 0.5150 1.5800 1.0550 0.6200 1.0550
                 0.6200 0.6350 0.7400 0.6350 0.7400 0.9350 1.4600 0.9350 1.4600 0.3950 2.4200 0.3950 ;
    END
END OAI32XL

MACRO OAI32X4
    CLASS CORE ;
    FOREIGN OAI32X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1550 0.8200 4.2750 1.1500 ;
        RECT  2.3100 0.8200 4.2750 0.9400 ;
        RECT  1.8950 0.9700 2.4300 1.0900 ;
        RECT  2.0450 0.9400 2.4300 1.0900 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8450 1.1400 8.2150 1.3800 ;
        RECT  6.7550 1.0600 8.0550 1.1800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3500 1.2700 5.3150 1.3900 ;
        RECT  3.3500 1.0600 3.4700 1.3900 ;
        RECT  2.5550 1.0600 3.4700 1.1800 ;
        RECT  1.0150 1.2100 2.6750 1.3300 ;
        RECT  2.5550 1.0600 2.6750 1.3300 ;
        RECT  1.1750 1.2100 1.4350 1.3800 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4800 1.1750 8.6300 1.4350 ;
        RECT  6.1750 1.5000 8.6000 1.6200 ;
        RECT  8.4350 1.2400 8.6000 1.6200 ;
        RECT  7.3750 1.3000 7.6150 1.6200 ;
        RECT  6.1750 1.2200 6.2950 1.6200 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 1.5100 5.6550 1.6300 ;
        RECT  5.5350 1.2400 5.6550 1.6300 ;
        RECT  2.9900 1.3000 3.2300 1.6300 ;
        RECT  0.7350 1.2300 0.8550 1.6300 ;
        RECT  0.5950 1.2300 0.8550 1.3800 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8150 0.6500 9.0550 0.7700 ;
        RECT  6.2950 0.7600 8.9350 0.8800 ;
        RECT  7.9750 0.6500 8.2150 0.8800 ;
        RECT  7.9350 1.7400 8.0550 2.2100 ;
        RECT  1.8750 1.7500 8.0550 1.8700 ;
        RECT  7.1350 0.6500 7.3750 0.8800 ;
        RECT  6.6550 1.7400 6.7750 2.2100 ;
        RECT  6.2950 0.6500 6.5350 0.8800 ;
        RECT  5.9350 0.8200 6.4150 0.9400 ;
        RECT  5.8150 1.7500 6.0750 1.9600 ;
        RECT  5.9350 0.8200 6.0550 1.9600 ;
        RECT  4.4350 1.7500 4.5550 2.2100 ;
        RECT  1.8750 1.7500 1.9950 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  5.3950 0.3400 5.6350 0.4600 ;
        RECT  5.3950 -0.1800 5.5150 0.4600 ;
        RECT  4.4350 0.3400 4.6750 0.4600 ;
        RECT  4.4350 -0.1800 4.5550 0.4600 ;
        RECT  3.4750 0.3400 3.7150 0.4600 ;
        RECT  3.4750 -0.1800 3.5950 0.4600 ;
        RECT  2.5150 0.3400 2.7550 0.4600 ;
        RECT  2.5150 -0.1800 2.6350 0.4600 ;
        RECT  1.5550 0.3400 1.7950 0.4600 ;
        RECT  1.5550 -0.1800 1.6750 0.4600 ;
        RECT  0.5950 0.3400 0.8350 0.4600 ;
        RECT  0.5950 -0.1800 0.7150 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.5750 1.7400 8.6950 2.7900 ;
        RECT  7.2350 1.9900 7.4750 2.1500 ;
        RECT  7.2350 1.9900 7.3550 2.7900 ;
        RECT  5.8150 2.0800 6.0550 2.2000 ;
        RECT  5.8150 2.0800 5.9350 2.7900 ;
        RECT  3.2700 1.9900 3.5100 2.1500 ;
        RECT  3.2700 1.9900 3.3900 2.7900 ;
        RECT  0.5950 1.7500 0.7150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.4150 0.6500 9.2950 0.6500 9.2950 0.5300 8.5750 0.5300 8.5750 0.6400 8.4550 0.6400
                 8.4550 0.5300 7.7350 0.5300 7.7350 0.6400 7.6150 0.6400 7.6150 0.5300 6.8950 0.5300
                 6.8950 0.6400 6.7750 0.6400 6.7750 0.5300 6.0550 0.5300 6.0550 0.7000 0.1150 0.7000
                 0.1150 0.5800 5.9350 0.5800 5.9350 0.4100 6.7750 0.4100 6.7750 0.4000 6.8950 0.4000
                 6.8950 0.4100 7.6150 0.4100 7.6150 0.4000 7.7350 0.4000 7.7350 0.4100 8.4550 0.4100
                 8.4550 0.4000 8.5750 0.4000 8.5750 0.4100 9.4150 0.4100 ;
    END
END OAI32X4

MACRO OAI32X2
    CLASS CORE ;
    FOREIGN OAI32X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0350 1.0600 4.5350 1.1800 ;
        RECT  3.2600 1.0600 3.4100 1.4350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5550 0.8200 2.6750 1.1500 ;
        RECT  2.3900 0.8200 2.6750 1.1450 ;
        RECT  0.5950 0.8200 2.6750 0.9400 ;
        RECT  0.5950 0.8200 0.7150 1.1500 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5300 1.3000 3.7700 1.4200 ;
        RECT  3.5500 1.3000 3.7000 1.7250 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0600 2.2700 1.3000 ;
        RECT  2.1000 1.0600 2.2500 1.4350 ;
        RECT  0.9750 1.0600 2.2700 1.1800 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.3000 1.5700 1.4200 ;
        RECT  1.2300 1.4650 1.3800 1.7250 ;
        RECT  1.2600 1.3000 1.3800 1.7250 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2150 0.6500 4.4550 0.7700 ;
        RECT  3.3750 0.7600 4.3350 0.8800 ;
        RECT  3.5750 1.8450 3.6950 2.2100 ;
        RECT  3.3750 0.6500 3.6150 0.8800 ;
        RECT  2.7950 1.8450 3.6950 1.9650 ;
        RECT  2.7950 0.8200 3.4950 0.9400 ;
        RECT  2.7950 0.8200 2.9150 1.9650 ;
        RECT  1.6700 1.5600 2.9150 1.6800 ;
        RECT  2.6250 1.5200 2.9150 1.6800 ;
        RECT  1.6700 1.5600 1.7900 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  2.4750 0.3400 2.7150 0.4600 ;
        RECT  2.4750 -0.1800 2.5950 0.4600 ;
        RECT  1.5150 0.3400 1.7550 0.4600 ;
        RECT  1.5150 -0.1800 1.6350 0.4600 ;
        RECT  0.5550 0.3400 0.7950 0.4600 ;
        RECT  0.5550 -0.1800 0.6750 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  4.2150 1.5600 4.3350 2.7900 ;
        RECT  2.8150 2.0850 3.0550 2.2050 ;
        RECT  2.8150 2.0850 2.9350 2.7900 ;
        RECT  0.5550 1.5600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8150 0.6500 4.6950 0.6500 4.6950 0.5300 3.9750 0.5300 3.9750 0.6400 3.8550 0.6400
                 3.8550 0.5300 3.1350 0.5300 3.1350 0.7000 0.0750 0.7000 0.0750 0.5800 3.0150 0.5800
                 3.0150 0.4100 3.8550 0.4100 3.8550 0.4000 3.9750 0.4000 3.9750 0.4100 4.8150 0.4100 ;
    END
END OAI32X2

MACRO OAI32X1
    CLASS CORE ;
    FOREIGN OAI32X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0750 0.8150 2.2500 1.2150 ;
        RECT  2.0750 0.8150 2.1950 1.2250 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 1.0500 1.1100 1.4750 ;
        RECT  0.9400 1.3550 1.0900 1.7600 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.3500 1.6700 1.7250 ;
        RECT  1.5350 1.2350 1.6550 1.7250 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.4500 0.8000 1.8700 ;
        RECT  0.6500 1.1350 0.7700 1.8700 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3300 1.0450 0.5100 1.4350 ;
        RECT  0.3300 1.0350 0.4500 1.4350 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4268  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2700 0.9950 1.9350 1.1150 ;
        RECT  1.8150 0.6450 1.9350 1.1150 ;
        RECT  1.2700 0.9950 1.3900 2.2050 ;
        RECT  1.2300 1.1750 1.3900 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  0.9150 0.5150 1.1550 0.6350 ;
        RECT  0.9150 -0.1800 1.0350 0.6350 ;
        RECT  0.1350 -0.1800 0.2550 0.6950 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  2.0350 1.5550 2.1550 2.7900 ;
        RECT  0.1700 1.5550 0.2900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3550 0.6950 2.2350 0.6950 2.2350 0.5250 1.5150 0.5250 1.5150 0.8750 0.5550 0.8750
                 0.5550 0.6350 0.6750 0.6350 0.6750 0.7550 1.3950 0.7550 1.3950 0.4050 2.3550 0.4050 ;
    END
END OAI32X1

MACRO OAI31XL
    CLASS CORE ;
    FOREIGN OAI31XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.1250 1.3800 1.6150 ;
        RECT  1.2300 1.1250 1.3800 1.5850 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 0.8850 1.7000 1.2700 ;
        RECT  1.5800 0.8750 1.7000 1.2700 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.8850 0.5100 1.3400 ;
        RECT  0.3600 0.8850 0.4800 1.3650 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.3350 1.0900 1.7250 ;
        RECT  0.9400 1.1450 1.0600 1.7250 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6000 1.4650 1.9600 1.7250 ;
        RECT  1.8400 0.5250 1.9600 1.7250 ;
        RECT  1.4200 1.7350 1.7200 1.8550 ;
        RECT  1.6000 1.4650 1.7200 1.8550 ;
        RECT  1.4200 1.7350 1.5400 1.9750 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.0000 -0.1800 1.1200 0.7650 ;
        RECT  0.1600 -0.1800 0.2800 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.8400 1.8450 1.9600 2.7900 ;
        RECT  0.4600 1.8450 0.5800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6000 0.7050 1.4000 0.7050 1.4000 1.0050 0.6300 1.0050 0.6300 0.7650 0.5800 0.7650
                 0.5800 0.5250 0.7000 0.5250 0.7000 0.6450 0.7500 0.6450 0.7500 0.8850 1.2800 0.8850
                 1.2800 0.5850 1.6000 0.5850 ;
    END
END OAI31XL

MACRO OAI31X4
    CLASS CORE ;
    FOREIGN OAI31X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7900 0.9700 4.2950 1.0900 ;
        RECT  3.7900 0.8200 3.9100 1.0900 ;
        RECT  2.2000 0.8200 3.9100 0.9400 ;
        RECT  1.8550 0.9700 2.3200 1.0900 ;
        RECT  2.0450 0.9400 2.3200 1.0900 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0950 1.0900 5.2150 1.3300 ;
        RECT  5.0000 0.8850 5.1500 1.2100 ;
        RECT  4.5650 1.0900 5.2150 1.2100 ;
        RECT  3.3400 1.2100 4.6850 1.3300 ;
        RECT  3.3400 1.0600 3.4600 1.3300 ;
        RECT  2.5450 1.0600 3.4600 1.1800 ;
        RECT  1.5250 1.2100 2.6650 1.3300 ;
        RECT  2.5450 1.0600 2.6650 1.3300 ;
        RECT  1.5250 0.9900 1.6450 1.3300 ;
        RECT  0.8750 0.9900 1.6450 1.1100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9300 1.4500 5.5550 1.5700 ;
        RECT  5.4350 1.2400 5.5550 1.5700 ;
        RECT  2.7850 1.3000 3.0250 1.5700 ;
        RECT  0.9300 1.3200 1.0500 1.5700 ;
        RECT  0.5950 1.3200 1.0500 1.4400 ;
        RECT  0.5950 1.2300 0.8550 1.4400 ;
        RECT  0.5950 1.2000 0.7150 1.4400 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3750 1.2250 7.0750 1.3450 ;
        RECT  6.6850 1.2250 6.9450 1.3800 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1072  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0950 0.6500 7.3350 0.7700 ;
        RECT  6.1350 0.7600 7.2150 0.8800 ;
        RECT  6.9150 1.5600 7.0350 2.2100 ;
        RECT  1.8350 1.6900 7.0350 1.8100 ;
        RECT  6.1350 0.6500 6.4950 0.8800 ;
        RECT  6.1350 1.4650 6.3100 1.8100 ;
        RECT  6.1350 0.6500 6.2550 1.8100 ;
        RECT  6.0750 1.5600 6.1950 2.2100 ;
        RECT  4.3950 1.6900 4.5150 2.2100 ;
        RECT  1.8350 1.6900 1.9550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  5.3550 0.3400 5.5950 0.4600 ;
        RECT  5.3550 -0.1800 5.4750 0.4600 ;
        RECT  4.3950 0.3400 4.6350 0.4600 ;
        RECT  4.3950 -0.1800 4.5150 0.4600 ;
        RECT  3.4350 0.3400 3.6750 0.4600 ;
        RECT  3.4350 -0.1800 3.5550 0.4600 ;
        RECT  2.4750 0.3400 2.7150 0.4600 ;
        RECT  2.4750 -0.1800 2.5950 0.4600 ;
        RECT  1.5150 0.3400 1.7550 0.4600 ;
        RECT  1.5150 -0.1800 1.6350 0.4600 ;
        RECT  0.5550 0.3400 0.7950 0.4600 ;
        RECT  0.5550 -0.1800 0.6750 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  7.3350 1.5600 7.4550 2.7900 ;
        RECT  6.4950 1.9300 6.6150 2.7900 ;
        RECT  5.6550 1.9300 5.7750 2.7900 ;
        RECT  3.0150 1.9300 3.1350 2.7900 ;
        RECT  0.4550 1.5600 0.5750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.6950 0.6500 7.5750 0.6500 7.5750 0.5300 6.8550 0.5300 6.8550 0.6400 6.7350 0.6400
                 6.7350 0.5300 6.0150 0.5300 6.0150 0.7000 0.0750 0.7000 0.0750 0.5800 5.8950 0.5800
                 5.8950 0.4100 6.7350 0.4100 6.7350 0.4000 6.8550 0.4000 6.8550 0.4100 7.6950 0.4100 ;
    END
END OAI31X4

MACRO OAI31X2
    CLASS CORE ;
    FOREIGN OAI31X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 0.9750 3.7000 1.4400 ;
        RECT  3.5500 0.9450 3.6700 1.4400 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6100 0.8850 2.8300 1.1450 ;
        RECT  0.6500 0.8200 2.8000 0.9400 ;
        RECT  2.6100 0.8200 2.7300 1.1500 ;
        RECT  0.6500 0.8200 0.7700 1.1500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9300 1.0600 2.4500 1.1800 ;
        RECT  1.2300 1.0600 1.3800 1.4350 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8700 1.3000 2.1100 1.4200 ;
        RECT  1.7550 1.5200 2.0150 1.6700 ;
        RECT  1.8700 1.3000 2.0150 1.6700 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5536  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3100 0.6500 3.6700 0.7700 ;
        RECT  1.7900 1.7900 3.4300 1.9100 ;
        RECT  3.3100 0.6500 3.4300 1.9100 ;
        RECT  2.9700 1.5600 3.4300 1.9100 ;
        RECT  3.1700 1.5600 3.2900 2.2100 ;
        RECT  2.9700 1.4650 3.1200 1.9100 ;
        RECT  1.7900 1.7900 1.9100 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  2.5300 0.3400 2.7700 0.4600 ;
        RECT  2.5300 -0.1800 2.6500 0.4600 ;
        RECT  1.5700 0.3400 1.8100 0.4600 ;
        RECT  1.5700 -0.1800 1.6900 0.4600 ;
        RECT  0.6100 0.3400 0.8500 0.4600 ;
        RECT  0.6100 -0.1800 0.7300 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.5900 1.5600 3.7100 2.7900 ;
        RECT  2.6900 2.0300 2.9300 2.1500 ;
        RECT  2.6900 2.0300 2.8100 2.7900 ;
        RECT  0.5100 1.5600 0.6300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.0300 0.6500 3.9100 0.6500 3.9100 0.5300 3.1900 0.5300 3.1900 0.7000 0.1300 0.7000
                 0.1300 0.5800 3.0700 0.5800 3.0700 0.4100 4.0300 0.4100 ;
    END
END OAI31X2

MACRO OAI31X1
    CLASS CORE ;
    FOREIGN OAI31X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.0300 1.3800 1.4850 ;
        RECT  1.2300 1.0000 1.3500 1.4850 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.0300 1.6700 1.4850 ;
        RECT  1.5500 1.0000 1.6700 1.4850 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.9850 0.4400 1.2450 ;
        RECT  0.3200 0.7600 0.4400 1.2450 ;
        RECT  0.0700 0.9850 0.2200 1.4400 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.0650 1.0900 1.4350 ;
        RECT  0.8400 1.0100 0.9600 1.3850 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3284  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3200 1.6050 1.9600 1.7250 ;
        RECT  1.8400 0.5900 1.9600 1.7250 ;
        RECT  1.8100 0.8850 1.9600 1.1450 ;
        RECT  1.3200 1.6050 1.4400 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.0000 -0.1800 1.1200 0.6400 ;
        RECT  0.1600 -0.1800 0.2800 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.7400 1.8450 1.8600 2.7900 ;
        RECT  0.3600 1.5600 0.4800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5400 0.8800 0.5800 0.8800 0.5800 0.5900 0.7000 0.5900 0.7000 0.7600 1.4200 0.7600
                 1.4200 0.5900 1.5400 0.5900 ;
    END
END OAI31X1

MACRO OAI2BB2XL
    CLASS CORE ;
    FOREIGN OAI2BB2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8000 0.8000 1.1450 ;
        RECT  0.6100 1.0000 0.7300 1.3450 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9700 1.0400 1.0900 1.5250 ;
        RECT  0.9400 1.0400 1.0900 1.4950 ;
        END
    END A0N
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.1300 2.8300 1.6000 ;
        RECT  2.6800 1.1000 2.8000 1.6000 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.1100 3.4100 1.4350 ;
        RECT  3.1900 1.2800 3.3100 1.6000 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1920  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9500 0.8900 3.0700 1.8400 ;
        RECT  2.9200 0.6800 3.0400 1.0100 ;
        RECT  2.6250 1.7200 3.0700 1.8400 ;
        RECT  2.4400 1.8400 2.8850 1.9600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  1.9600 -0.1800 2.0800 0.9200 ;
        RECT  0.6100 -0.1800 0.7300 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.0800 1.9600 3.3200 2.0800 ;
        RECT  3.0800 1.9600 3.2000 2.7900 ;
        RECT  1.8600 1.9000 1.9800 2.7900 ;
        RECT  0.7900 1.6450 0.9100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.4600 0.9200 3.3400 0.9200 3.3400 0.5600 2.6800 0.5600 2.6800 0.8000 2.6200 0.8000
                 2.6200 0.9200 2.5600 0.9200 2.5600 1.4000 1.4800 1.4000 1.4800 0.6800 1.6000 0.6800
                 1.6000 1.2800 2.4400 1.2800 2.4400 0.8000 2.5000 0.8000 2.5000 0.6800 2.5600 0.6800
                 2.5600 0.4400 3.4600 0.4400 ;
        POLYGON  2.4400 0.5200 2.3200 0.5200 2.3200 1.1600 1.7200 1.1600 1.7200 0.5600 0.9700 0.5600
                 0.9700 0.6800 0.2550 0.6800 0.2550 1.5250 0.4900 1.5250 0.4900 1.7650 0.3700 1.7650
                 0.3700 1.6450 0.1350 1.6450 0.1350 0.5600 0.8500 0.5600 0.8500 0.4400 1.8400 0.4400
                 1.8400 1.0400 2.2000 1.0400 2.2000 0.4000 2.4400 0.4000 ;
        POLYGON  1.8600 1.6400 1.3300 1.6400 1.3300 1.7650 1.2100 1.7650 1.2100 0.9200 1.0900 0.9200
                 1.0900 0.6800 1.2100 0.6800 1.2100 0.8000 1.3300 0.8000 1.3300 1.5200 1.8600 1.5200 ;
    END
END OAI2BB2XL

MACRO OAI2BB2X4
    CLASS CORE ;
    FOREIGN OAI2BB2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0100 0.5100 1.4650 ;
        RECT  0.3750 1.0100 0.4950 1.4950 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0200 0.8350 1.4000 ;
        RECT  0.6500 1.0650 0.8000 1.4350 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0250 1.2800 8.2650 1.4000 ;
        RECT  8.0250 1.2800 8.1450 1.5900 ;
        RECT  5.5750 1.4700 8.1450 1.5900 ;
        RECT  6.5550 1.3000 6.7950 1.5900 ;
        RECT  5.5250 1.5200 5.7850 1.6700 ;
        RECT  5.5750 1.2800 5.6950 1.6700 ;
        RECT  5.4250 1.2800 5.6950 1.4000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.1740  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.4028  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8150 0.9400 6.0750 1.1700 ;
        RECT  5.8450 0.9400 5.9650 1.3500 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9650 0.4600 8.2050 0.5800 ;
        RECT  6.3750 0.4100 8.0850 0.5300 ;
        RECT  5.9850 1.7100 7.7850 1.8300 ;
        RECT  7.1250 0.4100 7.3650 0.5800 ;
        RECT  6.2250 0.4600 6.5250 0.5800 ;
        RECT  5.1850 0.7000 6.3450 0.8200 ;
        RECT  6.2250 0.4600 6.3450 0.8200 ;
        RECT  5.9850 1.7100 6.1050 2.0100 ;
        RECT  5.1850 1.7900 6.1050 1.9100 ;
        RECT  5.4450 0.6500 5.6850 0.8200 ;
        RECT  2.6450 1.6900 5.3050 1.8100 ;
        RECT  5.1850 0.7000 5.3050 1.9100 ;
        RECT  4.9450 1.5200 5.3050 1.8100 ;
        RECT  4.1250 1.5600 4.2450 2.0100 ;
        RECT  2.6450 1.6900 2.7650 2.0100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  4.5450 -0.1800 4.7850 0.3400 ;
        RECT  3.6450 0.4600 3.8850 0.5800 ;
        RECT  3.6450 -0.1800 3.7650 0.5800 ;
        RECT  2.8050 0.4600 3.0450 0.5800 ;
        RECT  2.8050 -0.1800 2.9250 0.5800 ;
        RECT  2.0250 -0.1800 2.1450 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  8.2450 2.1900 8.4850 2.3100 ;
        RECT  8.2450 2.1900 8.3650 2.7900 ;
        RECT  6.7550 2.1900 6.9950 2.3100 ;
        RECT  6.7550 2.1900 6.8750 2.7900 ;
        RECT  5.0850 2.2700 5.3250 2.7900 ;
        RECT  3.2850 2.1700 3.5250 2.2900 ;
        RECT  3.2850 2.1700 3.4050 2.7900 ;
        RECT  2.0050 1.9300 2.1250 2.7900 ;
        RECT  0.5550 1.6150 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.5650 0.8300 8.5050 0.8300 8.5050 2.0700 6.6350 2.0700 6.6350 2.2500 5.7200 2.2500
                 5.7200 2.1500 4.7800 2.1500 4.7800 2.2500 3.6450 2.2500 3.6450 2.0500 3.1600 2.0500
                 3.1600 2.2500 2.2450 2.2500 2.2450 1.8100 1.3050 1.8100 1.3050 1.0800 1.4250 1.0800
                 1.4250 0.6500 1.6650 0.6500 1.6650 0.7700 1.5450 0.7700 1.5450 1.0800 2.0250 1.0800
                 2.0250 1.2100 2.5050 1.2100 2.5050 0.8300 2.4450 0.8300 2.4450 0.5900 2.5650 0.5900
                 2.5650 0.7000 3.2850 0.7000 3.2850 0.5900 3.4050 0.5900 3.4050 0.7000 4.1250 0.7000
                 4.1250 0.5900 4.2450 0.5900 4.2450 0.7000 4.8800 0.7000 4.8800 0.4600 5.2050 0.4600
                 5.2050 0.4100 5.9850 0.4100 5.9850 0.4600 6.1050 0.4600 6.1050 0.5800 5.8650 0.5800
                 5.8650 0.5300 5.3250 0.5300 5.3250 0.5800 5.0000 0.5800 5.0000 0.8200 4.2450 0.8200
                 4.2450 0.8300 4.1250 0.8300 4.1250 0.8200 3.4050 0.8200 3.4050 0.8300 3.2850 0.8300
                 3.2850 0.8200 2.6250 0.8200 2.6250 1.3300 1.9050 1.3300 1.9050 1.2000 1.4250 1.2000
                 1.4250 1.6900 2.3650 1.6900 2.3650 2.1300 3.0400 2.1300 3.0400 1.9300 3.7650 1.9300
                 3.7650 2.1300 4.6600 2.1300 4.6600 2.0300 5.8400 2.0300 5.8400 2.1300 6.5150 2.1300
                 6.5150 1.9500 8.3850 1.9500 8.3850 0.8300 6.8250 0.8300 6.8250 0.7700 6.7050 0.7700
                 6.7050 0.6500 6.9450 0.6500 6.9450 0.7100 7.5450 0.7100 7.5450 0.6500 7.7850 0.6500
                 7.7850 0.7100 8.4450 0.7100 8.4450 0.5900 8.5650 0.5900 ;
        POLYGON  7.5350 1.1800 6.4350 1.1800 6.4350 1.2900 6.1950 1.2900 6.1950 1.1700 6.3150 1.1700
                 6.3150 1.0600 7.5350 1.0600 ;
        POLYGON  5.0050 1.4000 3.3250 1.4000 3.3250 1.5700 1.6650 1.5700 1.6650 1.4400 1.5450 1.4400
                 1.5450 1.3200 1.7850 1.3200 1.7850 1.4500 3.0850 1.4500 3.0850 1.2800 5.0050 1.2800 ;
        RECT  2.7450 1.0000 4.0250 1.1200 ;
        POLYGON  2.3850 1.0900 2.1450 1.0900 2.1450 0.9600 1.7850 0.9600 1.7850 0.4800 0.9150 0.4800
                 0.9150 0.8900 0.2400 0.8900 0.2400 1.5850 0.2550 1.5850 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.7050 0.1200 1.7050 0.1200 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000
                 0.2550 0.7700 0.7950 0.7700 0.7950 0.3600 1.9050 0.3600 1.9050 0.8400 2.2650 0.8400
                 2.2650 0.9700 2.3850 0.9700 ;
        POLYGON  1.1850 1.2500 1.1550 1.2500 1.1550 1.6800 1.0950 1.6800 1.0950 2.2100 0.9750 2.2100
                 0.9750 1.5600 1.0350 1.5600 1.0350 0.6000 1.1550 0.6000 1.1550 1.0100 1.1850 1.0100 ;
    END
END OAI2BB2X4

MACRO OAI2BB2X2
    CLASS CORE ;
    FOREIGN OAI2BB2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.1850 0.5650 1.4000 ;
        RECT  0.3550 1.1850 0.4750 1.5950 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.5200 0.8550 1.7150 ;
        RECT  0.7350 1.3100 0.8550 1.7150 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.5250 4.8650 1.6450 ;
        RECT  4.7450 1.2200 4.8650 1.6450 ;
        RECT  3.5850 1.2300 4.0450 1.3800 ;
        RECT  3.7850 1.2300 3.9050 1.6450 ;
        RECT  3.5850 1.2300 3.9050 1.4200 ;
        RECT  3.5850 1.1800 3.7050 1.4200 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3650 1.1800 4.6250 1.4050 ;
        RECT  4.1650 1.2000 4.6250 1.4000 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.5250 0.6500 4.7650 0.7700 ;
        RECT  3.3450 0.9400 4.6450 1.0600 ;
        RECT  4.5250 0.6500 4.6450 1.0600 ;
        RECT  4.0650 1.7650 4.1850 2.2100 ;
        RECT  3.3450 1.7650 4.1850 1.8850 ;
        RECT  3.6850 0.6500 3.9250 0.7700 ;
        RECT  3.6850 0.6500 3.8050 1.0600 ;
        RECT  3.3450 0.9400 3.4650 1.8850 ;
        RECT  2.3350 1.5500 3.4650 1.6700 ;
        RECT  2.5450 1.5500 2.6650 2.2100 ;
        RECT  2.3350 1.5200 2.5950 1.6700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  2.8450 0.4600 3.0850 0.5800 ;
        RECT  2.8450 -0.1800 2.9650 0.5800 ;
        RECT  2.0050 0.4600 2.2450 0.5800 ;
        RECT  2.0050 -0.1800 2.1250 0.5800 ;
        RECT  0.6150 -0.1800 0.7350 0.8250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.7050 1.7650 4.8250 2.7900 ;
        RECT  3.2650 2.0050 3.5050 2.1500 ;
        RECT  3.2650 2.0050 3.3850 2.7900 ;
        RECT  1.9050 1.5600 2.0250 2.7900 ;
        RECT  0.5950 1.8350 0.7150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.1250 0.6500 5.0050 0.6500 5.0050 0.5300 4.2850 0.5300 4.2850 0.6500 4.1650 0.6500
                 4.1650 0.5300 3.4450 0.5300 3.4450 0.6500 3.4150 0.6500 3.4150 0.8200 1.7050 0.8200
                 1.7050 0.7700 1.5850 0.7700 1.5850 0.6500 1.8250 0.6500 1.8250 0.7000 2.4250 0.7000
                 2.4250 0.6500 2.6650 0.6500 2.6650 0.7000 3.2950 0.7000 3.2950 0.4100 5.1250 0.4100 ;
        POLYGON  3.2250 1.4000 1.2150 1.4000 1.2150 1.5200 1.1350 1.5200 1.1350 1.9550 1.0150 1.9550
                 1.0150 1.4000 1.0950 1.4000 1.0950 0.6000 1.2150 0.6000 1.2150 1.2800 3.2250 1.2800 ;
        POLYGON  2.4450 1.0900 1.3450 1.0900 1.3450 0.4800 0.9750 0.4800 0.9750 1.0650 0.1850 1.0650
                 0.1850 1.7150 0.2950 1.7150 0.2950 1.9550 0.1750 1.9550 0.1750 1.8350 0.0650 1.8350
                 0.0650 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000 0.2550 0.9450 0.8550 0.9450
                 0.8550 0.3600 1.4650 0.3600 1.4650 0.9700 2.4450 0.9700 ;
    END
END OAI2BB2X2

MACRO OAI2BB2X1
    CLASS CORE ;
    FOREIGN OAI2BB2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4450 1.1800 0.5650 1.6700 ;
        RECT  0.3050 1.1800 0.5650 1.4000 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.5200 1.1450 1.7050 ;
        RECT  0.8850 1.3300 1.0050 1.7050 ;
        END
    END A0N
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.1500 3.1200 1.4350 ;
        RECT  2.8550 1.1000 2.9750 1.3700 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 0.8850 3.7000 1.2000 ;
        RECT  3.4800 1.0800 3.6000 1.3900 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4750 1.5550 3.3600 1.6750 ;
        RECT  3.2400 0.8000 3.3600 1.6750 ;
        RECT  3.0950 0.8000 3.3600 0.9200 ;
        RECT  3.0950 0.6800 3.2150 0.9200 ;
        RECT  2.6750 1.5300 2.7950 2.1800 ;
        RECT  2.3350 1.5300 2.7950 1.6700 ;
        RECT  2.3350 1.5200 2.5950 1.6700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  2.1950 0.5500 2.4350 0.6700 ;
        RECT  2.1950 -0.1800 2.3150 0.6700 ;
        RECT  0.6850 -0.1800 0.8050 0.8200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.4800 1.5300 3.6000 2.7900 ;
        RECT  2.0350 1.5300 2.1550 2.7900 ;
        RECT  0.6250 1.8250 0.7450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.6350 0.7300 3.5150 0.7300 3.5150 0.6100 3.3850 0.6100 3.3850 0.5600 2.9750 0.5600
                 2.9750 0.9100 1.8350 0.9100 1.8350 0.6700 1.9550 0.6700 1.9550 0.7900 2.6150 0.7900
                 2.6150 0.7400 2.8550 0.7400 2.8550 0.4400 3.5050 0.4400 3.5050 0.4900 3.6350 0.4900 ;
        POLYGON  2.6950 1.2000 2.4550 1.2000 2.4550 1.1500 1.5950 1.1500 1.5950 0.4800 1.0450 0.4800
                 1.0450 1.0600 0.1850 1.0600 0.1850 1.7050 0.3250 1.7050 0.3250 1.9450 0.2050 1.9450
                 0.2050 1.8250 0.0650 1.8250 0.0650 0.7200 0.2050 0.7200 0.2050 0.6000 0.3250 0.6000
                 0.3250 0.9400 0.9250 0.9400 0.9250 0.3600 1.7150 0.3600 1.7150 1.0300 2.5750 1.0300
                 2.5750 1.0800 2.6950 1.0800 ;
        POLYGON  2.1550 1.3900 1.3850 1.3900 1.3850 1.9450 1.1650 1.9450 1.1650 2.0650 1.0450 2.0650
                 1.0450 1.8250 1.2650 1.8250 1.2650 0.8400 1.1650 0.8400 1.1650 0.6000 1.2850 0.6000
                 1.2850 0.7200 1.3850 0.7200 1.3850 1.2700 2.1550 1.2700 ;
    END
END OAI2BB2X1

MACRO OAI2BB1XL
    CLASS CORE ;
    FOREIGN OAI2BB1XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 0.8850 1.6700 1.3550 ;
        RECT  1.5500 0.8550 1.6700 1.3550 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.1600 1.5300 ;
        RECT  1.0400 1.1700 1.1600 1.5300 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1350 0.8000 1.5900 ;
        RECT  0.6800 1.1100 0.8000 1.5900 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4950 1.7100 0.6150 1.9500 ;
        RECT  0.4100 1.1100 0.5300 1.8300 ;
        RECT  0.1150 1.1100 0.5300 1.2300 ;
        RECT  0.1150 0.6300 0.3950 0.7500 ;
        RECT  0.2750 0.4900 0.3950 0.7500 ;
        RECT  0.0700 0.8850 0.2350 1.1450 ;
        RECT  0.1150 0.6300 0.2350 1.2300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  0.9150 -0.1800 1.0350 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.7750 2.2300 1.8950 2.7900 ;
        RECT  0.9750 2.2300 1.0950 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6750 0.7350 1.4000 0.7350 1.4000 1.4750 1.4550 1.4750 1.4550 1.8300 1.3350 1.8300
                 1.3350 1.5950 1.2800 1.5950 1.2800 0.9900 0.3550 0.9900 0.3550 0.8700 1.2800 0.8700
                 1.2800 0.6150 1.5550 0.6150 1.5550 0.4900 1.6750 0.4900 ;
    END
END OAI2BB1XL

MACRO OAI2BB1X4
    CLASS CORE ;
    FOREIGN OAI2BB1X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7950 1.0750 3.3750 1.1950 ;
        RECT  0.6800 1.0400 2.9150 1.1600 ;
        RECT  1.9150 1.0400 2.1550 1.1950 ;
        RECT  0.6500 1.0750 0.8000 1.4350 ;
        RECT  0.4350 1.0750 0.8000 1.1950 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4200 1.1750 4.5700 1.4350 ;
        RECT  4.1950 1.1750 4.5700 1.3150 ;
        RECT  4.1950 1.0750 4.3150 1.3150 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5950 1.0450 3.8350 1.1950 ;
        RECT  3.4950 0.9400 3.7550 1.1200 ;
        END
    END A0N
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1072  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0750 1.5550 3.1950 2.2100 ;
        RECT  0.0700 1.5550 3.1950 1.6750 ;
        RECT  2.3950 0.7350 2.6350 0.8550 ;
        RECT  0.1950 0.7850 2.5150 0.9050 ;
        RECT  2.2350 1.5550 2.3550 2.2100 ;
        RECT  1.3950 1.5550 1.5150 2.2100 ;
        RECT  0.9150 0.7350 1.1550 0.9050 ;
        RECT  0.5550 1.5550 0.6750 2.2100 ;
        RECT  0.1950 0.7850 0.3150 1.6750 ;
        RECT  0.0700 1.4650 0.2200 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  3.4950 -0.1800 3.6150 0.7250 ;
        RECT  1.6550 0.5450 1.8950 0.6650 ;
        RECT  1.6550 -0.1800 1.7750 0.6650 ;
        RECT  0.2750 0.5450 0.5150 0.6650 ;
        RECT  0.2750 -0.1800 0.3950 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  4.3350 1.5600 4.4550 2.7900 ;
        RECT  3.4950 1.5600 3.6150 2.7900 ;
        RECT  2.6550 1.7950 2.7750 2.7900 ;
        RECT  1.8150 1.7950 1.9350 2.7900 ;
        RECT  0.9750 1.7950 1.0950 2.7900 ;
        RECT  0.1350 1.8450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.2550 0.9550 4.0750 0.9550 4.0750 1.5550 4.0350 1.5550 4.0350 2.2100 3.9150 2.2100
                 3.9150 1.4350 1.2950 1.4350 1.2950 1.4000 1.1750 1.4000 1.1750 1.2800 1.4150 1.2800
                 1.4150 1.3150 2.4350 1.3150 2.4350 1.2800 2.6750 1.2800 2.6750 1.3150 3.9550 1.3150
                 3.9550 0.8350 4.1350 0.8350 4.1350 0.6750 4.2550 0.6750 ;
    END
END OAI2BB1X4

MACRO OAI2BB1X2
    CLASS CORE ;
    FOREIGN OAI2BB1X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.1750 2.8300 1.4350 ;
        RECT  2.5150 1.1750 2.8300 1.2950 ;
        RECT  2.5150 1.0550 2.6350 1.2950 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 1.0000 2.1550 1.1500 ;
        RECT  1.7550 0.9400 2.0150 1.1200 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4350 1.0400 1.6350 1.1600 ;
        RECT  0.6500 1.0400 0.8000 1.4350 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5536  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.5550 1.5150 2.2100 ;
        RECT  0.0700 1.5550 1.5150 1.6750 ;
        RECT  0.1950 0.8000 1.0950 0.9200 ;
        RECT  0.9750 0.6300 1.0950 0.9200 ;
        RECT  0.5550 1.5550 0.6750 2.2100 ;
        RECT  0.1950 0.8000 0.3150 1.6750 ;
        RECT  0.0700 1.4650 0.2200 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.6150 -0.1800 1.7350 0.6800 ;
        RECT  0.3350 -0.1800 0.4550 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.6450 2.2000 2.7650 2.7900 ;
        RECT  1.8750 2.2000 1.9950 2.7900 ;
        RECT  0.9750 1.7950 1.0950 2.7900 ;
        RECT  0.1350 1.8450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.6350 0.8100 2.3950 0.8100 2.3950 1.5200 2.3550 1.5200 2.3550 1.8000 2.2350 1.8000
                 2.2350 1.4000 1.0750 1.4000 1.0750 1.2800 2.2750 1.2800 2.2750 0.6900 2.6350 0.6900 ;
    END
END OAI2BB1X2

MACRO OAI2BB1X1
    CLASS CORE ;
    FOREIGN OAI2BB1X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1200 1.9600 1.4350 ;
        RECT  1.7400 0.9600 1.8600 1.2700 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 1.0350 1.3800 1.4700 ;
        RECT  1.2100 1.0100 1.3300 1.4700 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1650 1.0900 1.4350 ;
        RECT  0.8150 1.1650 1.0900 1.2850 ;
        RECT  0.8150 1.0350 0.9350 1.2850 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3284  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.3000 0.6750 2.1900 ;
        RECT  0.2550 1.3000 0.6750 1.4200 ;
        RECT  0.2550 0.6000 0.3750 1.4200 ;
        RECT  0.0700 0.8850 0.3750 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.7750 2.2300 1.8950 2.7900 ;
        RECT  0.9750 1.5900 1.0950 2.7900 ;
        RECT  0.1350 1.5400 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.8100 0.8400 1.6200 0.8400 1.6200 1.7100 1.5150 1.7100 1.5150 1.8300 1.3950 1.8300
                 1.3950 1.5900 1.5000 1.5900 1.5000 0.8900 0.6150 0.8900 0.6150 1.1800 0.4950 1.1800
                 0.4950 0.7700 1.5000 0.7700 1.5000 0.7200 1.6900 0.7200 1.6900 0.6000 1.8100 0.6000 ;
    END
END OAI2BB1X1

MACRO OAI22XL
    CLASS CORE ;
    FOREIGN OAI22XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.3600 1.3800 1.7250 ;
        RECT  1.2100 1.2800 1.3300 1.6500 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1650 1.6700 1.6200 ;
        RECT  1.5300 1.1000 1.6500 1.6200 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0800 0.5100 1.5300 ;
        RECT  0.3600 1.0800 0.4800 1.5550 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.9800 0.8200 1.4050 ;
        RECT  0.6500 1.1750 0.8000 1.5850 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2172  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2800 0.8600 1.5800 0.9800 ;
        RECT  1.4600 0.6800 1.5800 0.9800 ;
        RECT  0.9700 1.0400 1.4000 1.1600 ;
        RECT  1.2800 0.8600 1.4000 1.1600 ;
        RECT  0.9700 1.0400 1.0900 1.8600 ;
        RECT  0.9400 1.4650 1.0900 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.6900 1.7400 1.8100 2.7900 ;
        RECT  0.2200 1.7400 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.0000 0.9200 1.8800 0.9200 1.8800 0.5600 1.1600 0.5600 1.1600 0.9200 1.0400 0.9200
                 1.0400 0.8600 0.0750 0.8600 0.0750 0.7400 1.0400 0.7400 1.0400 0.4400 2.0000 0.4400 ;
    END
END OAI22XL

MACRO OAI22X4
    CLASS CORE ;
    FOREIGN OAI22X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0550 1.0600 7.1750 1.1800 ;
        RECT  4.1300 1.0600 4.2800 1.4350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5350 0.9900 3.6950 1.1100 ;
        RECT  2.9150 0.9400 3.1750 1.1100 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6750 1.3000 6.1950 1.4200 ;
        RECT  4.6550 1.5200 4.9150 1.6700 ;
        RECT  4.6750 1.3000 4.9150 1.6700 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5150 1.2600 3.0350 1.3800 ;
        RECT  2.6250 1.2300 2.8850 1.3800 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8550 0.6500 7.0950 0.7700 ;
        RECT  4.3350 0.7600 6.9750 0.8800 ;
        RECT  6.0150 0.6500 6.2550 0.8800 ;
        RECT  5.8750 1.5600 5.9950 2.2100 ;
        RECT  1.7350 1.7900 5.9950 1.9100 ;
        RECT  5.1750 0.6500 5.4150 0.8800 ;
        RECT  4.5950 1.7900 4.7150 2.2100 ;
        RECT  4.3350 0.6500 4.5750 0.8800 ;
        RECT  3.8150 0.8200 4.4550 0.9400 ;
        RECT  3.7850 1.7900 4.0450 1.9600 ;
        RECT  3.8150 0.8200 3.9350 1.9600 ;
        RECT  3.1150 1.5600 3.2350 2.2100 ;
        RECT  1.7350 1.5600 1.8550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  3.4350 0.3400 3.6750 0.4600 ;
        RECT  3.4350 -0.1800 3.5550 0.4600 ;
        RECT  2.4750 0.3400 2.7150 0.4600 ;
        RECT  2.4750 -0.1800 2.5950 0.4600 ;
        RECT  1.5150 0.3400 1.7550 0.4600 ;
        RECT  1.5150 -0.1800 1.6350 0.4600 ;
        RECT  0.5550 0.3400 0.7950 0.4600 ;
        RECT  0.5550 -0.1800 0.6750 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  6.5150 1.5600 6.6350 2.7900 ;
        RECT  5.1750 2.0300 5.4150 2.1500 ;
        RECT  5.1750 2.0300 5.2950 2.7900 ;
        RECT  3.7950 2.0800 4.0350 2.2000 ;
        RECT  3.7950 2.0800 3.9150 2.7900 ;
        RECT  2.3150 2.0300 2.5550 2.1500 ;
        RECT  2.3150 2.0300 2.4350 2.7900 ;
        RECT  1.0950 1.5600 1.2150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.4550 0.6500 7.3350 0.6500 7.3350 0.5300 6.6150 0.5300 6.6150 0.6400 6.4950 0.6400
                 6.4950 0.5300 5.7750 0.5300 5.7750 0.6400 5.6550 0.6400 5.6550 0.5300 4.9350 0.5300
                 4.9350 0.6400 4.8150 0.6400 4.8150 0.5300 4.0950 0.5300 4.0950 0.7000 0.0750 0.7000
                 0.0750 0.5800 3.9750 0.5800 3.9750 0.4100 4.8150 0.4100 4.8150 0.4000 4.9350 0.4000
                 4.9350 0.4100 5.6550 0.4100 5.6550 0.4000 5.7750 0.4000 5.7750 0.4100 6.4950 0.4100
                 6.4950 0.4000 6.6150 0.4000 6.6150 0.4100 7.4550 0.4100 ;
    END
END OAI22X4

MACRO OAI22X2
    CLASS CORE ;
    FOREIGN OAI22X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0600 3.3150 1.1800 ;
        RECT  2.3900 1.0600 2.5400 1.4350 ;
        RECT  2.1150 1.1800 2.5400 1.3000 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6350 0.9700 1.7550 1.2100 ;
        RECT  1.4650 0.9400 1.7250 1.0900 ;
        RECT  0.4150 0.9700 1.7550 1.0900 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.4650 3.1200 1.7250 ;
        RECT  2.9700 1.3000 3.0900 1.7250 ;
        RECT  2.7350 1.3000 3.0900 1.4200 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.2800 1.1550 1.4000 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.2800 0.8000 1.7250 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0150 0.6500 3.2550 0.7700 ;
        RECT  2.1500 0.7600 3.1350 0.8800 ;
        RECT  2.6550 1.5550 2.7750 2.2100 ;
        RECT  1.1350 1.5550 2.7750 1.6750 ;
        RECT  2.1500 0.6500 2.4150 0.8800 ;
        RECT  1.8750 0.9400 2.2700 1.0600 ;
        RECT  2.1500 0.6500 2.2700 1.0600 ;
        RECT  1.7550 1.5200 2.0150 1.6750 ;
        RECT  1.8750 0.9400 1.9950 1.6750 ;
        RECT  1.1350 1.5550 1.2550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  1.3350 0.4600 1.5750 0.5800 ;
        RECT  1.3350 -0.1800 1.4550 0.5800 ;
        RECT  0.4950 0.4600 0.7350 0.5800 ;
        RECT  0.4950 -0.1800 0.6150 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.2950 1.5600 3.4150 2.7900 ;
        RECT  1.8550 1.7950 2.0950 2.1500 ;
        RECT  1.8550 1.7950 1.9750 2.7900 ;
        RECT  0.4950 1.8450 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.6150 0.6500 3.4950 0.6500 3.4950 0.5300 2.7750 0.5300 2.7750 0.6400 2.6550 0.6400
                 2.6550 0.5300 1.9350 0.5300 1.9350 0.8200 0.1950 0.8200 0.1950 0.7700 0.0750 0.7700
                 0.0750 0.6500 0.3150 0.6500 0.3150 0.7000 0.9150 0.7000 0.9150 0.6500 1.1550 0.6500
                 1.1550 0.7000 1.8150 0.7000 1.8150 0.4100 2.6550 0.4100 2.6550 0.4000 2.7750 0.4000
                 2.7750 0.4100 3.6150 0.4100 ;
    END
END OAI22X2

MACRO OAI22X1
    CLASS CORE ;
    FOREIGN OAI22X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.4100 1.3800 1.7250 ;
        RECT  1.2100 1.2400 1.3300 1.5350 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 0.9650 1.6700 1.4400 ;
        RECT  1.5200 0.9850 1.6700 1.4350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0600 0.5100 1.4350 ;
        RECT  0.2400 1.0500 0.4800 1.2400 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0850 0.8200 1.5000 ;
        RECT  0.7000 1.0700 0.8200 1.5000 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3489  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 0.7250 1.5150 0.8450 ;
        RECT  1.3950 0.6050 1.5150 0.8450 ;
        RECT  0.9700 1.0000 1.3350 1.1200 ;
        RECT  1.2150 0.7250 1.3350 1.1200 ;
        RECT  0.9700 1.0000 1.0900 2.2100 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  0.4950 0.5200 0.7350 0.6400 ;
        RECT  0.4950 -0.1800 0.6150 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.7100 1.5600 1.8300 2.7900 ;
        RECT  0.2200 1.5600 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 0.7000 1.8150 0.7000 1.8150 0.4850 1.0950 0.4850 1.0950 0.8800 0.1350 0.8800
                 0.1350 0.6400 0.2550 0.6400 0.2550 0.7600 0.9750 0.7600 0.9750 0.3650 1.9350 0.3650 ;
    END
END OAI22X1

MACRO OAI222XL
    CLASS CORE ;
    FOREIGN OAI222XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1400 1.9600 1.6100 ;
        END
    END B0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.1400 2.8300 1.6100 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1400 0.8850 1.4700 ;
        RECT  0.6500 1.1400 0.8000 1.4750 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1600 2.3750 1.2800 ;
        RECT  2.2550 1.0250 2.3750 1.2800 ;
        RECT  2.1000 1.1600 2.2500 1.4350 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1400 0.5100 1.5150 ;
        RECT  0.3900 0.9600 0.5100 1.5150 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5150 1.1500 1.6700 1.6100 ;
        RECT  1.5150 1.1400 1.6350 1.6100 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4116  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2550 1.7300 3.0700 1.8500 ;
        RECT  2.9500 0.9000 3.0700 1.8500 ;
        RECT  2.6350 0.9000 3.0700 1.0200 ;
        RECT  2.7350 1.7300 2.8550 2.0900 ;
        RECT  2.6350 0.7200 2.7550 1.0200 ;
        RECT  2.6800 1.7300 2.8550 2.0150 ;
        RECT  2.5150 0.6000 2.6350 0.8400 ;
        RECT  1.2550 1.7300 1.3750 2.0900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  0.9850 -0.1800 1.1050 0.4500 ;
        RECT  0.1350 -0.1800 0.2550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.0950 1.9700 2.2150 2.7900 ;
        RECT  0.2850 1.9700 0.4050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1150 0.7800 2.8750 0.7800 2.8750 0.4800 2.2150 0.4800 2.2150 0.8400 2.0950 0.8400
                 2.0950 0.4800 1.4350 0.4800 1.4350 0.7800 1.1950 0.7800 1.1950 0.6600 1.3150 0.6600
                 1.3150 0.3600 2.9950 0.3600 2.9950 0.6600 3.1150 0.6600 ;
        POLYGON  1.7950 1.0200 0.6300 1.0200 0.6300 0.8400 0.4450 0.8400 0.4450 0.7200 0.7500 0.7200
                 0.7500 0.9000 1.6750 0.9000 1.6750 0.6000 1.7950 0.6000 ;
    END
END OAI222XL

MACRO OAI222X4
    CLASS CORE ;
    FOREIGN OAI222X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9600 1.0600 6.3600 1.1800 ;
        RECT  4.9450 1.2300 5.2050 1.3800 ;
        RECT  4.9600 1.0600 5.2050 1.3800 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 1.0600 9.5600 1.3000 ;
        RECT  9.2950 1.0600 9.5550 1.3800 ;
        RECT  8.1000 1.0600 9.5600 1.1800 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3100 1.0600 2.8300 1.1800 ;
        RECT  1.4650 1.0600 1.7250 1.3800 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0300 1.1750 7.1800 1.4350 ;
        RECT  4.1800 1.5000 7.1500 1.6200 ;
        RECT  7.0300 1.1750 7.1500 1.6200 ;
        RECT  5.3250 1.3000 5.5650 1.6200 ;
        RECT  4.1800 1.2200 4.3000 1.6200 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6100 1.5000 9.8800 1.6200 ;
        RECT  9.7600 1.2200 9.8800 1.6200 ;
        RECT  8.7200 1.3000 8.9600 1.6200 ;
        RECT  7.6100 1.1750 7.7600 1.6200 ;
        RECT  7.4600 1.2800 7.7600 1.4000 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5700 1.5000 3.4100 1.6200 ;
        RECT  3.2600 1.1750 3.4100 1.6200 ;
        RECT  1.9700 1.3000 2.2100 1.6200 ;
        RECT  0.5700 1.2800 0.6900 1.6200 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.7984  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.2200 1.4650 10.3700 1.7250 ;
        RECT  1.5300 1.7400 10.3400 1.8600 ;
        RECT  10.2200 0.6500 10.3400 1.8600 ;
        RECT  7.7000 0.8200 10.3400 0.9400 ;
        RECT  9.3800 0.6500 9.5000 0.9400 ;
        RECT  9.2800 1.7400 9.4000 2.2100 ;
        RECT  8.5400 0.6500 8.6600 0.9400 ;
        RECT  8.0000 1.7400 8.1200 2.2100 ;
        RECT  7.7000 0.6500 7.8200 0.9400 ;
        RECT  6.4400 1.7400 6.5600 2.2100 ;
        RECT  4.7600 1.7400 4.8800 2.2100 ;
        RECT  2.8100 1.7400 2.9300 2.2100 ;
        RECT  1.5300 1.7400 1.6500 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  3.5300 -0.1800 3.6500 0.7000 ;
        RECT  2.6900 -0.1800 2.8100 0.7000 ;
        RECT  1.8500 -0.1800 1.9700 0.7000 ;
        RECT  1.0100 -0.1800 1.1300 0.7000 ;
        RECT  0.1700 -0.1800 0.2900 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  9.8600 1.9800 10.1000 2.1500 ;
        RECT  9.8600 1.9800 9.9800 2.7900 ;
        RECT  8.5800 1.9800 8.8200 2.1500 ;
        RECT  8.5800 1.9800 8.7000 2.7900 ;
        RECT  7.2200 1.9800 7.4600 2.1500 ;
        RECT  7.2200 1.9800 7.3400 2.7900 ;
        RECT  5.6050 1.9800 5.8450 2.1500 ;
        RECT  5.6050 1.9800 5.7250 2.7900 ;
        RECT  3.8600 1.9800 4.1000 2.1500 ;
        RECT  3.8600 1.9800 3.9800 2.7900 ;
        RECT  2.1100 1.9800 2.3500 2.1500 ;
        RECT  2.1100 1.9800 2.2300 2.7900 ;
        RECT  0.8900 1.7400 1.0100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.7600 0.7000 10.6400 0.7000 10.6400 0.5300 9.9200 0.5300 9.9200 0.7000 9.8000 0.7000
                 9.8000 0.5300 9.0800 0.5300 9.0800 0.7000 8.9600 0.7000 8.9600 0.5300 8.2400 0.5300
                 8.2400 0.7000 8.1200 0.7000 8.1200 0.5300 7.4000 0.5300 7.4000 0.7000 7.2800 0.7000
                 7.2800 0.5300 6.5600 0.5300 6.5600 0.7000 6.4400 0.7000 6.4400 0.5300 5.7200 0.5300
                 5.7200 0.7000 5.6000 0.7000 5.6000 0.5300 4.8800 0.5300 4.8800 0.7000 4.7600 0.7000
                 4.7600 0.5300 4.0400 0.5300 4.0400 0.7000 3.9200 0.7000 3.9200 0.4100 10.7600 0.4100 ;
        POLYGON  6.9800 0.9400 0.5900 0.9400 0.5900 0.6500 0.7100 0.6500 0.7100 0.8200 1.4300 0.8200
                 1.4300 0.6500 1.5500 0.6500 1.5500 0.8200 2.2700 0.8200 2.2700 0.6500 2.3900 0.6500
                 2.3900 0.8200 3.1100 0.8200 3.1100 0.6500 3.2300 0.6500 3.2300 0.8200 4.3400 0.8200
                 4.3400 0.6500 4.4600 0.6500 4.4600 0.8200 5.1800 0.8200 5.1800 0.6500 5.3000 0.6500
                 5.3000 0.8200 6.0200 0.8200 6.0200 0.6500 6.1400 0.6500 6.1400 0.8200 6.8600 0.8200
                 6.8600 0.6500 6.9800 0.6500 ;
    END
END OAI222X4

MACRO OAI222X2
    CLASS CORE ;
    FOREIGN OAI222X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1500 1.1550 3.4650 1.3800 ;
        RECT  2.9700 1.1550 3.4650 1.3550 ;
        END
    END B1
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.5050 1.0100 4.6250 1.4200 ;
        RECT  4.3650 1.1500 4.6250 1.3800 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1650 1.2150 1.3800 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 1.2250 5.4450 1.3450 ;
        RECT  5.0000 1.1750 5.1500 1.4350 ;
        RECT  4.0850 1.5400 5.1200 1.6600 ;
        RECT  5.0000 1.1750 5.1200 1.6600 ;
        RECT  4.0850 1.2200 4.2050 1.6600 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.5000 3.7850 1.6200 ;
        RECT  3.6650 1.2200 3.7850 1.6200 ;
        RECT  2.6800 1.1750 2.8300 1.6200 ;
        RECT  2.4450 1.2800 2.8300 1.4000 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5350 1.5000 1.7150 1.6200 ;
        RECT  1.5200 1.2200 1.7150 1.6200 ;
        RECT  1.5200 1.1750 1.6700 1.6200 ;
        RECT  0.5350 1.2200 0.6550 1.6200 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.8992  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5650 1.4650 5.7300 1.7250 ;
        RECT  1.1150 1.7800 5.6850 1.9000 ;
        RECT  5.5650 0.7700 5.6850 1.9000 ;
        RECT  4.3450 0.7700 5.6850 0.8900 ;
        RECT  5.1850 0.6000 5.3050 0.8900 ;
        RECT  4.5650 1.7800 4.6850 2.2100 ;
        RECT  4.3450 0.6000 4.4650 0.8900 ;
        RECT  2.9850 1.7400 3.1050 2.2100 ;
        RECT  1.1150 1.7400 1.2350 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  1.8550 -0.1800 1.9750 0.7300 ;
        RECT  1.0150 -0.1800 1.1350 0.7300 ;
        RECT  0.1750 -0.1800 0.2950 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1450 2.0200 5.3850 2.1500 ;
        RECT  5.1450 2.0200 5.2650 2.7900 ;
        RECT  3.8650 2.0200 4.1050 2.1500 ;
        RECT  3.8650 2.0200 3.9850 2.7900 ;
        RECT  2.1850 2.0200 2.4250 2.1500 ;
        RECT  2.1850 2.0200 2.3050 2.7900 ;
        RECT  0.3750 1.7400 0.4950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7250 0.6500 5.6050 0.6500 5.6050 0.4800 4.8850 0.4800 4.8850 0.6500 4.7650 0.6500
                 4.7650 0.4800 4.0450 0.4800 4.0450 0.6500 3.9250 0.6500 3.9250 0.4800 3.2050 0.4800
                 3.2050 0.6500 3.0850 0.6500 3.0850 0.4800 2.3650 0.4800 2.3650 0.6500 2.2450 0.6500
                 2.2450 0.3600 5.7250 0.3600 ;
        POLYGON  3.6250 0.9700 0.5950 0.9700 0.5950 0.6800 0.7150 0.6800 0.7150 0.8500 1.4350 0.8500
                 1.4350 0.6800 1.5550 0.6800 1.5550 0.8500 2.6650 0.8500 2.6650 0.6000 2.7850 0.6000
                 2.7850 0.8500 3.5050 0.8500 3.5050 0.6000 3.6250 0.6000 ;
    END
END OAI222X2

MACRO OAI222X1
    CLASS CORE ;
    FOREIGN OAI222X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0900 0.7850 2.2500 1.2150 ;
        RECT  2.0900 0.7700 2.2100 1.2150 ;
        END
    END B0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.0300 2.8500 1.4350 ;
        RECT  2.7300 1.0150 2.8500 1.4350 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1150 1.0900 1.4350 ;
        RECT  0.8600 1.0100 0.9800 1.3200 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.7700 2.5400 1.2200 ;
        RECT  2.4100 0.7700 2.5300 1.2600 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0400 0.5100 1.4950 ;
        RECT  0.3900 1.0100 0.5100 1.4950 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.0300 1.6900 1.4350 ;
        RECT  1.5700 1.0150 1.6900 1.4350 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7811  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.4650 3.1200 1.7250 ;
        RECT  2.9700 0.7750 3.0900 1.7250 ;
        RECT  2.8900 1.5550 3.0100 2.2100 ;
        RECT  2.6700 0.7750 3.0900 0.8950 ;
        RECT  1.4100 1.5550 3.1200 1.6750 ;
        RECT  2.6700 0.6000 2.7900 0.8950 ;
        RECT  1.4100 1.5550 1.5300 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  1.0200 -0.1800 1.1400 0.6500 ;
        RECT  0.1800 -0.1800 0.3000 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.2500 1.7950 2.3700 2.7900 ;
        RECT  0.3800 1.6150 0.5000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.2100 0.6500 3.0900 0.6500 3.0900 0.5300 2.9100 0.5300 2.9100 0.4800 2.3700 0.4800
                 2.3700 0.6500 2.2500 0.6500 2.2500 0.4800 1.5300 0.4800 1.5300 0.6500 1.4100 0.6500
                 1.4100 0.3600 3.0300 0.3600 3.0300 0.4100 3.2100 0.4100 ;
        POLYGON  1.9500 0.8900 0.6000 0.8900 0.6000 0.6000 0.7200 0.6000 0.7200 0.7700 1.8300 0.7700
                 1.8300 0.6000 1.9500 0.6000 ;
    END
END OAI222X1

MACRO OAI221XL
    CLASS CORE ;
    FOREIGN OAI221XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0650 2.2900 1.4350 ;
        RECT  2.1700 1.0600 2.2900 1.4350 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.9800 1.9600 1.4350 ;
        RECT  1.8100 0.9800 1.9300 1.4650 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7800 1.3650 0.9000 1.6350 ;
        RECT  0.6500 1.4650 0.8000 1.7500 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0400 1.2550 1.4350 1.4100 ;
        RECT  1.1100 1.2200 1.4350 1.4100 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1750 0.5100 1.5950 ;
        RECT  0.3600 0.9600 0.4800 1.5950 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3120  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5300 0.6800 2.6500 0.9200 ;
        RECT  2.3900 1.7550 2.5400 2.0150 ;
        RECT  2.2900 1.5850 2.5300 1.9450 ;
        RECT  2.4100 0.8000 2.5300 2.0150 ;
        RECT  1.0200 1.5850 2.5300 1.7050 ;
        RECT  1.0200 1.5850 1.1400 1.9450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.0000 -0.1800 1.1200 0.5300 ;
        RECT  0.1350 -0.1800 0.2550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.6600 1.8250 1.7800 2.7900 ;
        RECT  0.3000 1.8250 0.4200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2300 0.9200 2.1100 0.9200 2.1100 0.6200 1.4500 0.6200 1.4500 0.8600 1.2100 0.8600
                 1.2100 0.7400 1.3300 0.7400 1.3300 0.5000 2.2300 0.5000 ;
        POLYGON  1.8700 0.8600 1.6900 0.8600 1.6900 1.1000 0.6300 1.1000 0.6300 0.8400 0.4600 0.8400
                 0.4600 0.7200 0.7500 0.7200 0.7500 0.9800 1.5700 0.9800 1.5700 0.7400 1.8700 0.7400 ;
    END
END OAI221XL

MACRO OAI221X4
    CLASS CORE ;
    FOREIGN OAI221X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7300 1.2300 8.4300 1.3500 ;
        RECT  7.8450 1.2300 8.1050 1.3800 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1050 1.2300 6.3650 1.3800 ;
        RECT  6.1050 1.0600 6.3300 1.3800 ;
        RECT  4.9900 1.0600 6.3300 1.1800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1950 1.0100 2.9400 1.1300 ;
        RECT  1.1750 1.2300 1.4350 1.3800 ;
        RECT  1.1950 1.0100 1.4350 1.3800 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7400 1.1750 6.8900 1.4350 ;
        RECT  4.3100 1.5000 6.8600 1.6200 ;
        RECT  6.7400 1.1750 6.8600 1.6200 ;
        RECT  5.6800 1.3000 5.9200 1.6200 ;
        RECT  4.3100 1.2200 4.4300 1.6200 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.5000 3.5400 1.6200 ;
        RECT  3.4200 1.2400 3.5400 1.6200 ;
        RECT  2.0200 1.2500 2.1400 1.6200 ;
        RECT  0.6800 1.1750 0.8000 1.6200 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        RECT  0.5600 1.3000 0.8000 1.4200 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5232  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5500 0.8850 8.9200 1.1450 ;
        RECT  7.7300 0.7700 8.6900 0.8900 ;
        RECT  8.5700 0.6000 8.6900 1.1450 ;
        RECT  1.1200 1.7400 8.6700 1.8600 ;
        RECT  8.3700 1.5600 8.6700 1.8600 ;
        RECT  8.5500 0.7200 8.6700 1.8600 ;
        RECT  8.3700 1.5600 8.4900 2.2100 ;
        RECT  7.7300 0.6000 7.8500 0.8900 ;
        RECT  7.5300 1.5600 7.6500 2.2100 ;
        RECT  6.2400 1.7400 6.3600 2.2100 ;
        RECT  4.9600 1.7400 5.0800 2.2100 ;
        RECT  2.9200 1.7400 3.0400 2.2100 ;
        RECT  1.1200 1.7400 1.2400 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        RECT  3.5600 -0.1800 3.6800 0.6500 ;
        RECT  2.7200 -0.1800 2.8400 0.6500 ;
        RECT  1.8800 -0.1800 2.0000 0.6500 ;
        RECT  1.0400 -0.1800 1.1600 0.6500 ;
        RECT  0.2000 -0.1800 0.3200 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        RECT  8.7900 1.5600 8.9100 2.7900 ;
        RECT  7.8900 1.9800 8.1300 2.1500 ;
        RECT  7.8900 1.9800 8.0100 2.7900 ;
        RECT  7.0500 1.9800 7.2900 2.1500 ;
        RECT  7.0500 1.9800 7.1700 2.7900 ;
        RECT  5.5400 1.9800 5.7800 2.1500 ;
        RECT  5.5400 1.9800 5.6600 2.7900 ;
        RECT  3.5000 1.9800 3.7400 2.1500 ;
        RECT  3.5000 1.9800 3.6200 2.7900 ;
        RECT  1.7000 1.9800 1.9400 2.1500 ;
        RECT  1.7000 1.9800 1.8200 2.7900 ;
        RECT  0.4800 1.7400 0.6000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.1100 0.6500 8.9900 0.6500 8.9900 0.4800 8.2700 0.4800 8.2700 0.6500 8.1500 0.6500
                 8.1500 0.4800 7.4300 0.4800 7.4300 0.6500 7.3100 0.6500 7.3100 0.4800 6.5900 0.4800
                 6.5900 0.6500 6.4700 0.6500 6.4700 0.4800 5.7500 0.4800 5.7500 0.6500 5.6300 0.6500
                 5.6300 0.4800 4.9100 0.4800 4.9100 0.6500 4.7900 0.6500 4.7900 0.4800 4.0700 0.4800
                 4.0700 0.6500 3.9500 0.6500 3.9500 0.3600 9.1100 0.3600 ;
        POLYGON  7.0700 0.7800 6.9500 0.7800 6.9500 0.8900 0.6200 0.8900 0.6200 0.6000 0.7400 0.6000
                 0.7400 0.7700 1.4600 0.7700 1.4600 0.6000 1.5800 0.6000 1.5800 0.7700 2.3000 0.7700
                 2.3000 0.6000 2.4200 0.6000 2.4200 0.7700 3.1400 0.7700 3.1400 0.6000 3.2600 0.6000
                 3.2600 0.7700 4.3700 0.7700 4.3700 0.6000 4.4900 0.6000 4.4900 0.7700 5.2100 0.7700
                 5.2100 0.6000 5.3300 0.6000 5.3300 0.7700 6.0500 0.7700 6.0500 0.6000 6.1700 0.6000
                 6.1700 0.7700 6.8300 0.7700 6.8300 0.6600 7.0700 0.6600 ;
    END
END OAI221X4

MACRO OAI221X2
    CLASS CORE ;
    FOREIGN OAI221X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1600 0.8500 4.2800 1.4400 ;
        RECT  4.1300 0.8500 4.2800 1.3050 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0550 1.1400 3.2950 1.3300 ;
        RECT  2.9150 1.1650 3.1750 1.3800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.1650 1.4350 1.3800 ;
        RECT  1.0550 1.1600 1.2950 1.3500 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6750 1.5000 3.7600 1.6200 ;
        RECT  3.5500 1.2200 3.7600 1.6200 ;
        RECT  3.5500 1.1750 3.7000 1.6200 ;
        RECT  2.6750 1.2200 2.7950 1.6200 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.5000 1.6900 1.6200 ;
        RECT  1.5700 1.2200 1.6900 1.6200 ;
        RECT  0.6800 1.1750 0.8000 1.6200 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        RECT  0.5300 1.3000 0.8000 1.4200 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7616  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4000 1.1750 4.5700 1.4350 ;
        RECT  4.4200 0.6800 4.5400 0.9200 ;
        RECT  1.0900 1.7400 4.5200 1.8600 ;
        RECT  4.2200 1.5600 4.5200 1.8600 ;
        RECT  4.4000 0.8000 4.5200 1.8600 ;
        RECT  4.2200 1.5600 4.3400 2.2100 ;
        RECT  3.1600 1.7400 3.2800 2.2100 ;
        RECT  1.0900 1.7400 1.2100 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  1.9300 -0.1800 2.0500 0.7300 ;
        RECT  1.0900 -0.1800 1.2100 0.7300 ;
        RECT  0.2500 -0.1800 0.3700 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  4.6400 1.5600 4.7600 2.7900 ;
        RECT  3.7400 1.9800 3.9800 2.1500 ;
        RECT  3.7400 1.9800 3.8600 2.7900 ;
        RECT  1.6700 1.9800 1.9100 2.1500 ;
        RECT  1.6700 1.9800 1.7900 2.7900 ;
        RECT  0.4500 1.7400 0.5700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.9600 0.7300 4.8400 0.7300 4.8400 0.5600 4.1200 0.5600 4.1200 0.7300 4.0000 0.7300
                 4.0000 0.5600 3.2800 0.5600 3.2800 0.7300 3.1600 0.7300 3.1600 0.5600 2.4400 0.5600
                 2.4400 0.7300 2.3200 0.7300 2.3200 0.4400 4.9600 0.4400 ;
        POLYGON  3.7600 0.8600 3.6400 0.8600 3.6400 0.9700 0.6700 0.9700 0.6700 0.6800 0.7900 0.6800
                 0.7900 0.8500 1.5100 0.8500 1.5100 0.6800 1.6300 0.6800 1.6300 0.8500 2.7400 0.8500
                 2.7400 0.6800 2.8600 0.6800 2.8600 0.8500 3.5200 0.8500 3.5200 0.7400 3.7600 0.7400 ;
    END
END OAI221X2

MACRO OAI221X1
    CLASS CORE ;
    FOREIGN OAI221X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.9850 2.5400 1.4400 ;
        RECT  2.4050 0.8950 2.5250 1.4400 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8850 1.0000 2.0050 1.3500 ;
        RECT  1.8100 1.0850 1.9600 1.4350 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1400 1.0900 1.4350 ;
        RECT  0.8350 1.1000 0.9550 1.3800 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.0350 1.6700 1.4900 ;
        RECT  1.5450 1.0100 1.6650 1.4900 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0100 0.5100 1.4950 ;
        RECT  0.3600 1.0100 0.5100 1.4650 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7639  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3850 1.6100 2.7800 1.7300 ;
        RECT  2.6600 0.7450 2.7800 1.7300 ;
        RECT  2.6450 0.6000 2.7650 0.8650 ;
        RECT  2.4450 1.5600 2.7800 1.7300 ;
        RECT  2.4450 1.5600 2.5650 2.2100 ;
        RECT  2.3900 1.6100 2.5650 2.0150 ;
        RECT  1.3850 1.6100 1.5050 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  0.9950 -0.1800 1.1150 0.6500 ;
        RECT  0.1550 -0.1800 0.2750 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.0250 1.8500 2.1450 2.7900 ;
        RECT  0.3550 1.6150 0.4750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3450 0.6500 2.2250 0.6500 2.2250 0.5300 2.0450 0.5300 2.0450 0.4800 1.5050 0.4800
                 1.5050 0.6500 1.3850 0.6500 1.3850 0.3600 2.1650 0.3600 2.1650 0.4100 2.3450 0.4100 ;
        POLYGON  1.9250 0.8800 1.7650 0.8800 1.7650 0.8900 0.5750 0.8900 0.5750 0.6000 0.6950 0.6000
                 0.6950 0.7700 1.6450 0.7700 1.6450 0.7600 1.8050 0.7600 1.8050 0.6000 1.9250 0.6000 ;
    END
END OAI221X1

MACRO OAI21XL
    CLASS CORE ;
    FOREIGN OAI21XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.0400 1.3800 1.5100 ;
        RECT  1.2300 1.0400 1.3500 1.5400 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.4650 1.0250 1.6600 ;
        RECT  0.9050 1.4200 1.0250 1.6600 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.3250 0.5100 1.7800 ;
        RECT  0.3850 1.3000 0.5050 1.7800 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5000 1.4650 1.6700 1.7250 ;
        RECT  1.5000 0.8000 1.6200 1.7800 ;
        RECT  1.4850 0.6800 1.6050 0.9200 ;
        RECT  1.1450 1.6600 1.6200 1.7800 ;
        RECT  1.0650 1.7800 1.2650 1.9000 ;
        RECT  1.0650 1.7800 1.1850 2.0200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.6450 -0.1800 0.7650 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.4850 1.9000 1.6050 2.7900 ;
        RECT  0.4250 1.9000 0.5450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1850 0.9200 1.1100 0.9200 1.1100 1.1600 0.2250 1.1600 0.2250 0.6800 0.3450 0.6800
                 0.3450 1.0400 0.9900 1.0400 0.9900 0.8000 1.0650 0.8000 1.0650 0.6800 1.1850 0.6800 ;
    END
END OAI21XL

MACRO OAI21X4
    CLASS CORE ;
    FOREIGN OAI21X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0550 1.2300 4.7550 1.3500 ;
        RECT  4.0550 1.2300 4.3350 1.3800 ;
        RECT  4.0550 1.1950 4.1750 1.4350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.1750 3.4100 1.4350 ;
        RECT  3.2350 0.9900 3.3800 1.2300 ;
        RECT  0.6150 0.9900 3.3800 1.1100 ;
        RECT  1.7750 0.9900 2.0150 1.1600 ;
        RECT  0.4950 1.0200 0.7350 1.1400 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1950 1.2800 2.6550 1.4000 ;
        RECT  1.1750 1.2300 1.4350 1.3800 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1072  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7750 0.7000 5.0150 0.8200 ;
        RECT  3.8150 0.8100 4.8950 0.9300 ;
        RECT  4.6350 1.5550 4.7550 2.2100 ;
        RECT  1.3550 1.5550 4.7550 1.6750 ;
        RECT  3.8150 0.7000 4.1750 0.9300 ;
        RECT  3.7950 1.5550 3.9900 2.0150 ;
        RECT  3.8150 0.7000 3.9350 2.0150 ;
        RECT  3.7950 1.5550 3.9150 2.2100 ;
        RECT  2.6350 1.5550 2.7550 2.2100 ;
        RECT  1.3550 1.5550 1.4750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  3.0950 0.5100 3.3350 0.6300 ;
        RECT  3.0950 -0.1800 3.2150 0.6300 ;
        RECT  2.2550 0.5100 2.4950 0.6300 ;
        RECT  2.2550 -0.1800 2.3750 0.6300 ;
        RECT  1.4150 0.5100 1.6550 0.6300 ;
        RECT  1.4150 -0.1800 1.5350 0.6300 ;
        RECT  0.5750 0.5100 0.8150 0.6300 ;
        RECT  0.5750 -0.1800 0.6950 0.6300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  5.0550 1.5600 5.1750 2.7900 ;
        RECT  4.2150 1.7950 4.3350 2.7900 ;
        RECT  3.3750 1.7950 3.4950 2.7900 ;
        RECT  1.9950 1.7950 2.1150 2.7900 ;
        RECT  0.4150 1.5600 0.5350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.3750 0.7000 5.2550 0.7000 5.2550 0.5800 4.5350 0.5800 4.5350 0.6900 4.4150 0.6900
                 4.4150 0.5800 3.6950 0.5800 3.6950 0.8700 0.2150 0.8700 0.2150 0.6300 0.3350 0.6300
                 0.3350 0.7500 1.0550 0.7500 1.0550 0.6300 1.1750 0.6300 1.1750 0.7500 1.8950 0.7500
                 1.8950 0.6300 2.0150 0.6300 2.0150 0.7500 2.7350 0.7500 2.7350 0.6300 2.8550 0.6300
                 2.8550 0.7500 3.5750 0.7500 3.5750 0.4600 4.4150 0.4600 4.4150 0.4500 4.5350 0.4500
                 4.5350 0.4600 5.3750 0.4600 ;
    END
END OAI21X4

MACRO OAI21X2
    CLASS CORE ;
    FOREIGN OAI21X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3600 1.0250 2.5400 1.4350 ;
        RECT  2.3600 1.0050 2.4800 1.4400 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1750 1.6700 1.4350 ;
        RECT  0.4800 1.0600 1.6400 1.1800 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.3000 1.0800 1.4200 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.3000 0.8000 1.7250 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5536  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1200 0.7650 2.4200 0.8850 ;
        RECT  2.3000 0.6450 2.4200 0.8850 ;
        RECT  1.0400 1.5550 2.2400 1.6750 ;
        RECT  2.1200 0.7650 2.2400 1.6750 ;
        RECT  2.1000 1.5550 2.2200 2.2100 ;
        RECT  1.8100 1.3150 2.2400 1.4350 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        RECT  1.0400 1.5550 1.1600 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  1.4600 -0.1800 1.5800 0.7000 ;
        RECT  0.6200 -0.1800 0.7400 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.5200 1.5600 2.6400 2.7900 ;
        RECT  1.6800 1.7950 1.8000 2.7900 ;
        RECT  0.4000 1.5600 0.5200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.8400 0.7000 2.7200 0.7000 2.7200 0.5250 2.0000 0.5250 2.0000 0.9400 0.2000 0.9400
                 0.2000 0.6500 0.3200 0.6500 0.3200 0.8200 1.0400 0.8200 1.0400 0.6500 1.1600 0.6500
                 1.1600 0.8200 1.8800 0.8200 1.8800 0.4050 2.8400 0.4050 ;
    END
END OAI21X2

MACRO OAI21X1
    CLASS CORE ;
    FOREIGN OAI21X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.0300 1.3800 1.4850 ;
        RECT  1.2300 1.0000 1.3500 1.4850 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.2000 1.0850 1.3200 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0000 0.5100 1.4850 ;
        RECT  0.3600 1.0000 0.5100 1.4550 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3284  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0650 1.6050 1.6700 1.7250 ;
        RECT  1.5000 1.4650 1.6700 1.7250 ;
        RECT  1.5000 0.7100 1.6200 1.7250 ;
        RECT  1.4850 0.5900 1.6050 0.8300 ;
        RECT  1.0650 1.6050 1.1850 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.6450 -0.1800 0.7650 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.4850 1.8450 1.6050 2.7900 ;
        RECT  0.4250 1.6050 0.5450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1850 0.8800 0.2250 0.8800 0.2250 0.5900 0.3450 0.5900 0.3450 0.7600 1.0650 0.7600
                 1.0650 0.5900 1.1850 0.5900 ;
    END
END OAI21X1

MACRO OAI211XL
    CLASS CORE ;
    FOREIGN OAI211XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3100 1.2500 1.4800 1.4900 ;
        RECT  1.2300 1.1750 1.4300 1.4350 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 1.1700 1.1100 1.5950 ;
        RECT  0.9400 1.1700 1.1100 1.5800 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.8000 1.6300 ;
        RECT  0.6700 1.1700 0.7900 1.6500 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.4650 0.5100 1.8650 ;
        RECT  0.3500 1.1700 0.4700 1.5850 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6000 1.7100 1.8950 1.9500 ;
        RECT  1.6150 0.5700 1.7350 0.8100 ;
        RECT  1.6000 0.6900 1.7200 1.9500 ;
        RECT  1.5200 1.7550 1.6700 2.0150 ;
        RECT  0.7700 1.7700 1.8950 1.8900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  0.5550 -0.1800 0.6750 0.8100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.3100 2.2300 1.4300 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1550 0.7500 1.0350 0.7500 1.0350 1.0500 0.1950 1.0500 0.1950 0.7500 0.0750 0.7500
                 0.0750 0.6300 0.3150 0.6300 0.3150 0.9300 0.9150 0.9300 0.9150 0.6300 1.1550 0.6300 ;
    END
END OAI211XL

MACRO OAI211X4
    CLASS CORE ;
    FOREIGN OAI211X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3050 1.2600 5.0850 1.3800 ;
        RECT  4.3650 1.2300 4.6250 1.3800 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0650 1.2000 6.7050 1.3200 ;
        RECT  6.5850 1.0800 6.7050 1.3200 ;
        RECT  6.4500 1.1750 6.6000 1.4350 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1950 1.0400 3.4350 1.1600 ;
        RECT  0.6800 0.9900 3.3150 1.1100 ;
        RECT  1.8350 0.9900 2.0750 1.1600 ;
        RECT  0.6500 1.0200 0.8000 1.4350 ;
        RECT  0.4350 1.0200 0.8000 1.1400 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 1.2800 2.7150 1.4000 ;
        RECT  2.3350 1.2300 2.5950 1.4000 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5232  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8250 0.8100 6.9650 0.9300 ;
        RECT  6.8450 0.6400 6.9650 0.9300 ;
        RECT  6.6050 1.5550 6.7250 2.2100 ;
        RECT  1.4150 1.5550 6.7250 1.6750 ;
        RECT  5.8250 0.7600 6.1250 0.9300 ;
        RECT  6.0050 0.6400 6.1250 0.9300 ;
        RECT  4.0650 0.9900 5.9450 1.1100 ;
        RECT  5.8250 0.7600 5.9450 1.1100 ;
        RECT  5.7650 1.5550 5.8850 2.2100 ;
        RECT  4.9250 1.5550 5.0450 2.2100 ;
        RECT  4.0650 1.5200 4.3350 1.6750 ;
        RECT  4.0850 1.5200 4.2050 2.2100 ;
        RECT  4.0650 0.9900 4.1850 1.6750 ;
        RECT  2.6950 1.5550 2.8150 2.2100 ;
        RECT  1.4150 1.5550 1.5350 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  3.4550 0.5100 3.6950 0.6300 ;
        RECT  3.4550 -0.1800 3.5750 0.6300 ;
        RECT  2.6150 0.5100 2.8550 0.6300 ;
        RECT  2.6150 -0.1800 2.7350 0.6300 ;
        RECT  1.7750 0.5100 2.0150 0.6300 ;
        RECT  1.7750 -0.1800 1.8950 0.6300 ;
        RECT  0.9350 0.5100 1.1750 0.6300 ;
        RECT  0.9350 -0.1800 1.0550 0.6300 ;
        RECT  0.1550 -0.1800 0.2750 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  7.0250 1.5600 7.1450 2.7900 ;
        RECT  6.1850 1.7950 6.3050 2.7900 ;
        RECT  5.3450 1.7950 5.4650 2.7900 ;
        RECT  4.4450 1.7950 4.6850 2.1500 ;
        RECT  4.4450 1.7950 4.5650 2.7900 ;
        RECT  3.6650 1.7950 3.7850 2.7900 ;
        RECT  2.0550 1.7950 2.1750 2.7900 ;
        RECT  0.3550 1.5600 0.4750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.3850 0.6900 7.2650 0.6900 7.2650 0.5200 6.5450 0.5200 6.5450 0.6900 6.4250 0.6900
                 6.4250 0.5200 5.7050 0.5200 5.7050 0.6900 5.5850 0.6900 5.5850 0.5200 4.9250 0.5200
                 4.9250 0.6300 4.6850 0.6300 4.6850 0.5200 4.0850 0.5200 4.0850 0.6300 3.8450 0.6300
                 3.8450 0.5100 3.9650 0.5100 3.9650 0.4000 7.3850 0.4000 ;
        POLYGON  5.3450 0.8200 5.2250 0.8200 5.2250 0.8700 0.5750 0.8700 0.5750 0.6300 0.6950 0.6300
                 0.6950 0.7500 1.4150 0.7500 1.4150 0.6300 1.5350 0.6300 1.5350 0.7500 2.2550 0.7500
                 2.2550 0.6300 2.3750 0.6300 2.3750 0.7500 3.0950 0.7500 3.0950 0.6300 3.2150 0.6300
                 3.2150 0.7500 4.2650 0.7500 4.2650 0.7000 4.5050 0.7000 4.5050 0.7500 5.1050 0.7500
                 5.1050 0.7000 5.3450 0.7000 ;
    END
END OAI211X4

MACRO OAI211X2
    CLASS CORE ;
    FOREIGN OAI211X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 1.0650 3.7000 1.4350 ;
        RECT  3.5250 1.0100 3.6450 1.3850 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.1800 2.6250 1.4250 ;
        RECT  2.2750 1.1800 2.6250 1.4000 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0400 1.6550 1.1600 ;
        RECT  0.3900 1.0400 0.5600 1.2800 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.2800 0.9950 1.4000 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.2800 0.8000 1.7250 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7616  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2850 0.6500 3.6450 0.7700 ;
        RECT  2.0350 0.9400 3.4050 1.0600 ;
        RECT  3.2850 0.6500 3.4050 1.0600 ;
        RECT  2.8750 1.5450 2.9950 2.2100 ;
        RECT  1.3750 1.5450 2.9950 1.6650 ;
        RECT  2.0350 0.9400 2.1550 2.2100 ;
        RECT  1.8100 1.1750 2.1550 1.6650 ;
        RECT  0.9750 1.5600 1.4950 1.6800 ;
        RECT  0.9750 1.5600 1.0950 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  1.7550 0.4600 1.9950 0.5800 ;
        RECT  1.7550 -0.1800 1.8750 0.5800 ;
        RECT  0.9150 0.4600 1.1550 0.5800 ;
        RECT  0.9150 -0.1800 1.0350 0.5800 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.2950 1.5600 3.4150 2.7900 ;
        RECT  2.4550 1.7850 2.5750 2.7900 ;
        RECT  1.6150 1.7850 1.7350 2.7900 ;
        RECT  0.3350 1.5600 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.0050 0.6500 3.8850 0.6500 3.8850 0.5300 3.1650 0.5300 3.1650 0.6500 3.0450 0.6500
                 3.0450 0.5300 2.3850 0.5300 2.3850 0.5800 2.1450 0.5800 2.1450 0.4600 2.2650 0.4600
                 2.2650 0.4100 4.0050 0.4100 ;
        POLYGON  2.8050 0.7700 2.6850 0.7700 2.6850 0.8200 0.5550 0.8200 0.5550 0.5800 0.6750 0.5800
                 0.6750 0.7000 1.3950 0.7000 1.3950 0.5800 1.5150 0.5800 1.5150 0.7000 2.5650 0.7000
                 2.5650 0.6500 2.8050 0.6500 ;
    END
END OAI211X2

MACRO OAI211X1
    CLASS CORE ;
    FOREIGN OAI211X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2800 1.3000 1.5200 1.4200 ;
        RECT  1.2800 0.5950 1.4000 1.4200 ;
        RECT  1.2300 0.5950 1.4000 0.8550 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9200 1.1950 1.1600 1.4000 ;
        RECT  0.9400 1.0400 1.0900 1.4350 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0400 0.8000 1.4350 ;
        RECT  0.5600 1.1150 0.8000 1.3200 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.4000 1.4000 ;
        RECT  0.2800 1.1600 0.4000 1.4000 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5104  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7800 1.5550 1.7600 1.6750 ;
        RECT  1.6400 0.7500 1.7600 1.6750 ;
        RECT  1.6200 1.5550 1.7400 2.2100 ;
        RECT  1.6200 0.6300 1.7400 0.8700 ;
        RECT  1.5200 1.5550 1.7400 2.0150 ;
        RECT  0.7800 1.5550 0.9000 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  0.5600 -0.1800 0.6800 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.2000 1.7950 1.3200 2.7900 ;
        RECT  0.1400 1.5600 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1000 0.9200 0.1400 0.9200 0.1400 0.6300 0.2600 0.6300 0.2600 0.8000 0.9800 0.8000
                 0.9800 0.6300 1.1000 0.6300 ;
    END
END OAI211X1

MACRO OA22XL
    CLASS CORE ;
    FOREIGN OA22XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0400 1.0200 1.1600 1.3300 ;
        RECT  0.9400 1.1200 1.0900 1.4350 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.9800 0.5100 1.4350 ;
        RECT  0.3600 0.9800 0.4800 1.7400 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 1.0800 0.8200 1.5200 ;
        RECT  0.6500 1.0800 0.8200 1.5000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.2700 1.6700 1.7250 ;
        RECT  1.5350 1.2600 1.6550 1.7400 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.4650 2.7650 1.6050 ;
        RECT  2.6450 0.6800 2.7650 1.6050 ;
        RECT  1.9750 1.8000 2.5400 1.9200 ;
        RECT  2.3900 1.4650 2.5400 1.9200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  2.1650 -0.1800 2.2850 0.4000 ;
        RECT  0.6150 -0.1800 0.7350 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.6150 1.8600 1.7350 2.7900 ;
        RECT  0.3350 1.8600 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.0750 1.1600 1.7900 1.1600 1.7900 1.1400 1.4000 1.1400 1.4000 1.6750 1.1550 1.6750
                 1.1550 1.9200 0.9150 1.9200 0.9150 1.8000 1.0350 1.8000 1.0350 1.5550 1.2800 1.5550
                 1.2800 0.7800 1.3950 0.7800 1.3950 0.6600 1.5150 0.6600 1.5150 0.9000 1.4000 0.9000
                 1.4000 1.0200 1.9100 1.0200 1.9100 1.0400 2.0750 1.0400 ;
        POLYGON  1.9350 0.9000 1.8150 0.9000 1.8150 0.5400 1.0950 0.5400 1.0950 0.9000 0.9750 0.9000
                 0.9750 0.8400 0.0750 0.8400 0.0750 0.7200 0.9750 0.7200 0.9750 0.4200 1.9350 0.4200 ;
    END
END OA22XL

MACRO OA22X4
    CLASS CORE ;
    FOREIGN OA22X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.2350 1.2950 ;
        RECT  1.1150 1.0550 1.2350 1.2950 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0100 0.5100 1.4650 ;
        RECT  0.3800 1.0100 0.5000 1.4950 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0300 0.8200 1.4350 ;
        RECT  0.7000 1.0200 0.8200 1.4350 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.8100 1.3400 1.9300 1.7250 ;
        RECT  1.6000 1.3400 1.9300 1.4600 ;
        RECT  1.6000 1.2200 1.7200 1.4600 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4050 1.1750 3.7000 1.4350 ;
        RECT  2.6850 0.7400 3.5850 0.8600 ;
        RECT  3.4650 0.6200 3.5850 0.8600 ;
        RECT  2.0800 1.3200 3.5250 1.4400 ;
        RECT  3.4050 0.7400 3.5250 1.4400 ;
        RECT  2.9200 1.3200 3.0400 2.2100 ;
        RECT  2.5650 0.6900 2.8050 0.8100 ;
        RECT  2.0800 1.3200 2.2000 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.8850 -0.1800 4.0050 0.6800 ;
        RECT  2.9850 0.5000 3.2250 0.6200 ;
        RECT  2.9850 -0.1800 3.1050 0.6200 ;
        RECT  2.2050 -0.1800 2.3250 0.6800 ;
        RECT  0.5550 -0.1800 0.6750 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.3400 1.5600 3.4600 2.7900 ;
        RECT  2.5000 1.5600 2.6200 2.7900 ;
        RECT  1.6600 1.8450 1.7800 2.7900 ;
        RECT  0.2200 1.6150 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.2850 1.1500 3.0450 1.1500 3.0450 1.1000 2.5400 1.1000 2.5400 1.1300 2.3000 1.1300
                 2.3000 1.1000 1.4800 1.1000 1.4800 1.6750 1.0950 1.6750 1.0950 2.2100 0.9750 2.2100
                 0.9750 1.5550 1.3600 1.5550 1.3600 0.7200 1.3950 0.7200 1.3950 0.6000 1.5150 0.6000
                 1.5150 0.8400 1.4800 0.8400 1.4800 0.9800 3.1650 0.9800 3.1650 1.0300 3.2850 1.0300 ;
        POLYGON  1.9350 0.6500 1.8150 0.6500 1.8150 0.4800 1.0950 0.4800 1.0950 0.8900 0.1350 0.8900
                 0.1350 0.6000 0.2550 0.6000 0.2550 0.7700 0.9750 0.7700 0.9750 0.3600 1.9350 0.3600 ;
    END
END OA22X4

MACRO OA22X2
    CLASS CORE ;
    FOREIGN OA22X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0250 1.4200 1.1950 1.6600 ;
        RECT  0.9400 1.4650 1.1350 1.7250 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.2800 0.5100 1.7400 ;
        RECT  0.3800 1.2800 0.5000 1.7600 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 1.2800 0.8200 1.7150 ;
        RECT  0.6500 1.3100 0.8000 1.7250 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4600 1.9600 1.7250 ;
        RECT  1.5550 1.4600 1.9600 1.5800 ;
        RECT  1.5550 1.4200 1.6750 1.6650 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.6500 2.7450 0.7700 ;
        RECT  2.2150 1.0050 2.5400 1.1450 ;
        RECT  2.3900 0.6500 2.5400 1.1450 ;
        RECT  2.2150 1.0050 2.3350 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.9850 -0.1800 3.1050 0.6400 ;
        RECT  2.0850 -0.1800 2.2050 0.5300 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.6350 1.5600 2.7550 2.7900 ;
        RECT  1.7950 1.8450 1.9150 2.7900 ;
        RECT  0.2200 1.8800 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.0950 1.3000 1.4350 1.3000 1.4350 1.9650 0.9150 1.9650 0.9150 1.8450 1.3150 1.8450
                 1.3150 0.8000 1.3950 0.8000 1.3950 0.6800 1.5150 0.6800 1.5150 0.9200 1.4350 0.9200
                 1.4350 1.1800 2.0950 1.1800 ;
        POLYGON  1.9350 0.9200 1.8150 0.9200 1.8150 0.5600 1.0950 0.5600 1.0950 1.1600 0.1950 1.1600
                 0.1950 0.8600 0.0750 0.8600 0.0750 0.7400 0.3150 0.7400 0.3150 1.0400 0.9750 1.0400
                 0.9750 0.4400 1.9350 0.4400 ;
    END
END OA22X2

MACRO OA22X1
    CLASS CORE ;
    FOREIGN OA22X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.2550 1.2950 ;
        RECT  1.1350 1.0550 1.2550 1.2950 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1650 0.5100 1.6200 ;
        RECT  0.3800 1.1000 0.5000 1.6200 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0000 0.8200 1.4350 ;
        RECT  0.7000 0.9800 0.8200 1.4350 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.6150 1.4000 1.9300 1.5200 ;
        RECT  1.6150 1.2800 1.7350 1.5200 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4200 0.6500 2.8250 0.7700 ;
        RECT  2.4200 0.6500 2.5400 1.1450 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.2750 1.0050 2.3950 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  2.1650 -0.1800 2.2850 0.5300 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.8550 1.8450 1.9750 2.7900 ;
        RECT  0.2200 1.7400 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.1550 1.1800 1.8550 1.1800 1.8550 1.1600 1.4950 1.1600 1.4950 1.8000 0.9950 1.8000
                 0.9950 1.6800 1.3750 1.6800 1.3750 0.8000 1.4750 0.8000 1.4750 0.6800 1.5950 0.6800
                 1.5950 0.9200 1.4950 0.9200 1.4950 1.0400 1.9750 1.0400 1.9750 1.0600 2.1550 1.0600 ;
        POLYGON  2.0150 0.9200 1.8950 0.9200 1.8950 0.5600 1.1750 0.5600 1.1750 0.9200 1.0550 0.9200
                 1.0550 0.8600 0.0750 0.8600 0.0750 0.7400 1.0550 0.7400 1.0550 0.4400 2.0150 0.4400 ;
    END
END OA22X1

MACRO OA21XL
    CLASS CORE ;
    FOREIGN OA21XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.5950 1.3800 0.9900 ;
        RECT  1.2300 0.5950 1.3500 1.2400 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7700 1.0200 0.8900 1.3300 ;
        RECT  0.6500 1.1750 0.8000 1.4950 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0400 0.5100 1.4800 ;
        RECT  0.3900 0.9600 0.5100 1.4800 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1300 0.7400 2.5350 0.8600 ;
        RECT  2.1000 0.8850 2.2500 1.1450 ;
        RECT  2.1300 0.7400 2.2500 1.1450 ;
        RECT  1.8500 1.0050 2.2500 1.1250 ;
        RECT  1.8500 1.0050 1.9700 1.7200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8900 -0.1800 2.0100 0.4000 ;
        RECT  0.6150 -0.1800 0.7350 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.4300 1.6000 1.5500 2.7900 ;
        RECT  0.2900 1.6000 0.4100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6900 1.4000 1.6200 1.4000 1.6200 1.4800 1.1300 1.4800 1.1300 1.7200 1.0100 1.7200
                 1.0100 1.3600 1.5000 1.3600 1.5000 0.6600 1.6200 0.6600 1.6200 1.1600 1.6900 1.1600 ;
        POLYGON  1.1100 0.9000 0.9900 0.9000 0.9900 0.8400 0.0750 0.8400 0.0750 0.7200 0.9900 0.7200
                 0.9900 0.6600 1.1100 0.6600 ;
    END
END OA21XL

MACRO OA21X4
    CLASS CORE ;
    FOREIGN OA21X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1750 1.6700 1.4350 ;
        RECT  1.3050 1.1750 1.6700 1.3400 ;
        RECT  1.3050 1.1000 1.4250 1.3400 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1350 1.1450 1.3800 ;
        RECT  0.8250 1.0900 1.0650 1.3100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0900 0.5100 1.5750 ;
        RECT  0.3600 1.0900 0.5100 1.5450 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1350 1.1750 3.4100 1.4350 ;
        RECT  2.0300 1.3200 3.2550 1.4400 ;
        RECT  3.1350 0.7100 3.2550 1.4400 ;
        RECT  3.0950 0.5900 3.2150 0.8800 ;
        RECT  2.2550 0.7600 3.2550 0.8800 ;
        RECT  2.8700 1.3200 2.9900 2.2100 ;
        RECT  2.2550 0.5900 2.3750 0.8800 ;
        RECT  2.0300 1.3200 2.1500 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.5150 -0.1800 3.6350 0.6400 ;
        RECT  2.6750 -0.1800 2.7950 0.6400 ;
        RECT  1.7750 -0.1800 1.8950 0.5300 ;
        RECT  0.6250 -0.1800 0.7450 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.2900 1.5600 3.4100 2.7900 ;
        RECT  2.4500 1.5600 2.5700 2.7900 ;
        RECT  1.6100 1.7950 1.7300 2.7900 ;
        RECT  0.4050 1.6950 0.5250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0150 1.1900 1.9100 1.1900 1.9100 1.6750 1.1650 1.6750 1.1650 2.2100 1.0450 2.2100
                 1.0450 1.5550 1.7900 1.5550 1.7900 0.9800 1.4650 0.9800 1.4650 0.6800 1.5850 0.6800
                 1.5850 0.8600 1.9100 0.8600 1.9100 1.0700 3.0150 1.0700 ;
        POLYGON  1.1650 0.9700 0.2050 0.9700 0.2050 0.6800 0.3250 0.6800 0.3250 0.8500 1.0450 0.8500
                 1.0450 0.6800 1.1650 0.6800 ;
    END
END OA21X4

MACRO OA21X2
    CLASS CORE ;
    FOREIGN OA21X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.7700 1.3800 1.1450 ;
        RECT  1.2500 0.7700 1.3700 1.2600 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.9500 1.2950 ;
        RECT  0.8300 1.0550 0.9500 1.2950 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1250 0.5100 1.5600 ;
        RECT  0.3900 1.0800 0.5100 1.5600 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1300 0.6500 2.4300 0.7700 ;
        RECT  1.8900 1.0050 2.2500 1.1450 ;
        RECT  2.1300 0.6500 2.2500 1.1450 ;
        RECT  2.1000 0.8850 2.2500 1.1450 ;
        RECT  1.8900 1.0050 2.0100 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.6700 -0.1800 2.7900 0.6400 ;
        RECT  1.7700 -0.1800 1.8900 0.5300 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3100 1.5600 2.4300 2.7900 ;
        RECT  1.4700 1.6200 1.5900 2.7900 ;
        RECT  0.3500 1.6800 0.4700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.7700 1.4800 1.6200 1.4800 1.6200 1.5000 1.1900 1.5000 1.1900 1.5350 1.1100 1.5350
                 1.1100 1.8000 0.9900 1.8000 0.9900 1.4150 1.0700 1.4150 1.0700 1.3800 1.5000 1.3800
                 1.5000 0.6800 1.6200 0.6800 1.6200 1.2400 1.7700 1.2400 ;
        POLYGON  1.1100 0.9200 0.9900 0.9200 0.9900 0.8600 0.0750 0.8600 0.0750 0.7400 0.9900 0.7400
                 0.9900 0.6800 1.1100 0.6800 ;
    END
END OA21X2

MACRO OA21X1
    CLASS CORE ;
    FOREIGN OA21X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.7700 1.3800 1.1450 ;
        RECT  1.2300 0.7700 1.3500 1.2600 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.9500 1.2950 ;
        RECT  0.8300 1.0550 0.9500 1.2950 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1250 0.5100 1.5600 ;
        RECT  0.3900 1.0800 0.5100 1.5600 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1300 0.6500 2.4300 0.7700 ;
        RECT  1.9700 1.0050 2.2500 1.1450 ;
        RECT  2.1300 0.6500 2.2500 1.1450 ;
        RECT  2.1000 0.8850 2.2500 1.1450 ;
        RECT  1.9700 1.0050 2.0900 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.7700 -0.1800 1.8900 0.5300 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.5500 1.6200 1.6700 2.7900 ;
        RECT  0.3500 1.6800 0.4700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.8200 1.4800 1.6200 1.4800 1.6200 1.5000 1.1900 1.5000 1.1900 1.8000 1.0700 1.8000
                 1.0700 1.3800 1.5000 1.3800 1.5000 0.6800 1.6200 0.6800 1.6200 1.2400 1.8200 1.2400 ;
        POLYGON  1.1100 0.9200 0.9900 0.9200 0.9900 0.8600 0.0750 0.8600 0.0750 0.7400 0.9900 0.7400
                 0.9900 0.6800 1.1100 0.6800 ;
    END
END OA21X1

MACRO NOR4XL
    CLASS CORE ;
    FOREIGN NOR4XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.0600 1.8000 1.2200 ;
        RECT  1.5200 1.1000 1.6700 1.4350 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2800 1.0500 1.4000 1.4750 ;
        RECT  1.2300 1.1750 1.3800 1.5850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.0500 1.0900 1.5050 ;
        RECT  0.9600 1.0500 1.0800 1.5350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1300 0.6150 1.3000 ;
        RECT  0.2950 1.1800 0.5650 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2544  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9200 0.8100 2.0400 1.5850 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  0.7000 0.8100 2.0400 0.9300 ;
        RECT  1.7900 1.4650 1.9600 1.7050 ;
        RECT  1.5400 0.4500 1.6600 0.9300 ;
        RECT  0.7000 0.4500 0.8200 0.9300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.9600 -0.1800 2.0800 0.6900 ;
        RECT  1.1200 -0.1800 1.2400 0.6900 ;
        RECT  0.2800 -0.1800 0.4000 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  0.4800 1.5100 0.6000 2.7900 ;
        END
    END VDD
END NOR4XL

MACRO NOR4X8
    CLASS CORE ;
    FOREIGN NOR4X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6050 1.2050 10.9850 1.3250 ;
        RECT  9.5850 1.2300 9.8450 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4800 1.1750 8.6300 1.4350 ;
        RECT  8.4800 1.0700 8.6000 1.4350 ;
        RECT  6.6550 1.1900 8.6300 1.3100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7150 1.2050 5.0750 1.3250 ;
        RECT  3.7850 1.2050 4.0450 1.3800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.1900 2.0750 1.3100 ;
        RECT  1.9550 1.0700 2.0750 1.3100 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.1393  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.9250 1.4650 12.0450 2.2100 ;
        RECT  9.4050 1.5000 12.0450 1.6200 ;
        RECT  0.6150 0.7900 11.6250 0.9100 ;
        RECT  11.5050 0.6700 11.6250 0.9100 ;
        RECT  11.0850 1.4650 11.2400 1.7250 ;
        RECT  11.1050 0.7900 11.2250 1.7250 ;
        RECT  11.0850 1.4650 11.2050 2.0100 ;
        RECT  10.6050 0.7400 10.8450 0.9100 ;
        RECT  10.2450 1.4700 10.3650 2.0100 ;
        RECT  9.7450 0.7400 9.9850 0.9100 ;
        RECT  9.4050 1.5000 9.5250 2.0100 ;
        RECT  8.9050 0.7400 9.1450 0.9100 ;
        RECT  8.0550 0.7400 8.2950 0.9100 ;
        RECT  7.2150 0.7400 7.4550 0.9100 ;
        RECT  6.3750 0.7400 6.6150 0.9100 ;
        RECT  5.5350 0.7400 5.7750 0.9100 ;
        RECT  4.6950 0.7400 4.9350 0.9100 ;
        RECT  3.8550 0.7400 4.0950 0.9100 ;
        RECT  3.0150 0.7400 3.2550 0.9100 ;
        RECT  2.1750 0.7400 2.4150 0.9100 ;
        RECT  1.3350 0.7400 1.5750 0.9100 ;
        RECT  0.4950 0.7400 0.7350 0.8600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.9250 -0.1800 12.0450 0.6700 ;
        RECT  11.0850 -0.1800 11.2050 0.6700 ;
        RECT  10.2450 -0.1800 10.3650 0.6700 ;
        RECT  9.3850 -0.1800 9.5050 0.6650 ;
        RECT  8.5350 -0.1800 8.6550 0.6700 ;
        RECT  7.6950 -0.1800 7.8150 0.6700 ;
        RECT  6.8550 -0.1800 6.9750 0.6700 ;
        RECT  6.0150 -0.1800 6.1350 0.6700 ;
        RECT  5.1750 -0.1800 5.2950 0.6700 ;
        RECT  4.3350 -0.1800 4.4550 0.6700 ;
        RECT  3.4950 -0.1800 3.6150 0.6650 ;
        RECT  2.6550 -0.1800 2.7750 0.6700 ;
        RECT  1.8150 -0.1800 1.9350 0.6700 ;
        RECT  0.9750 -0.1800 1.0950 0.6700 ;
        RECT  0.1350 -0.1800 0.2550 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  2.6550 1.7950 2.7750 2.7900 ;
        RECT  1.8150 1.7950 1.9350 2.7900 ;
        RECT  0.9750 1.7950 1.0950 2.7900 ;
        RECT  0.1350 1.4650 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6250 2.2500 8.9850 2.2500 8.9850 1.6750 8.2650 1.6750 8.2650 2.0100 8.1450 2.0100
                 8.1450 1.6750 7.3950 1.6750 7.3950 2.0100 7.2750 2.0100 7.2750 1.6750 6.5550 1.6750
                 6.5550 2.0100 6.4350 2.0100 6.4350 1.4650 6.5550 1.4650 6.5550 1.5550 7.2750 1.5550
                 7.2750 1.4650 7.3950 1.4650 7.3950 1.5550 8.1450 1.5550 8.1450 1.4700 8.2650 1.4700
                 8.2650 1.5550 8.9850 1.5550 8.9850 1.4700 9.1050 1.4700 9.1050 2.1300 9.8250 2.1300
                 9.8250 1.7400 9.9450 1.7400 9.9450 2.1300 10.6650 2.1300 10.6650 1.7400 10.7850 1.7400
                 10.7850 2.1300 11.5050 2.1300 11.5050 1.7400 11.6250 1.7400 ;
        POLYGON  8.6850 2.2500 6.0150 2.2500 6.0150 1.6200 5.2950 1.6200 5.2950 2.0100 5.1750 2.0100
                 5.1750 1.6200 4.4550 1.6200 4.4550 2.0100 4.3350 2.0100 4.3350 1.6200 3.6150 1.6200
                 3.6150 2.0100 3.4950 2.0100 3.4950 1.4700 3.6150 1.4700 3.6150 1.5000 4.3350 1.5000
                 4.3350 1.4700 4.4550 1.4700 4.4550 1.5000 5.1750 1.5000 5.1750 1.4650 5.2950 1.4650
                 5.2950 1.5000 6.0150 1.5000 6.0150 1.4650 6.1350 1.4650 6.1350 2.1300 6.8550 2.1300
                 6.8550 1.7950 6.9750 1.7950 6.9750 2.1300 7.6950 2.1300 7.6950 1.7950 7.8150 1.7950
                 7.8150 2.1300 8.5650 2.1300 8.5650 1.7950 8.6850 1.7950 ;
        POLYGON  5.7150 2.2500 3.0750 2.2500 3.0750 1.6750 2.3550 1.6750 2.3550 2.2100 2.2350 2.2100
                 2.2350 1.6750 1.5150 1.6750 1.5150 2.2100 1.3950 2.2100 1.3950 1.6750 0.6750 1.6750
                 0.6750 2.2100 0.5550 2.2100 0.5550 1.4650 0.6750 1.4650 0.6750 1.5550 1.3950 1.5550
                 1.3950 1.4650 1.5150 1.4650 1.5150 1.5550 2.2350 1.5550 2.2350 1.4700 2.3550 1.4700
                 2.3550 1.5550 3.0750 1.5550 3.0750 1.4700 3.1950 1.4700 3.1950 2.1300 3.9150 2.1300
                 3.9150 1.7400 4.0350 1.7400 4.0350 2.1300 4.7550 2.1300 4.7550 1.7400 4.8750 1.7400
                 4.8750 2.1300 5.5950 2.1300 5.5950 1.7400 5.7150 1.7400 ;
    END
END NOR4X8

MACRO NOR4X6
    CLASS CORE ;
    FOREIGN NOR4X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.1100 1.1700 7.7800 1.2900 ;
        RECT  7.2650 1.1700 7.5250 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8700 1.1750 6.0200 1.4350 ;
        RECT  5.8700 1.1100 5.9900 1.4350 ;
        RECT  5.1100 1.1750 6.0200 1.2950 ;
        RECT  4.9900 1.1500 5.2300 1.2700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.8900 1.1500 3.5100 1.2700 ;
        RECT  2.9150 1.1500 3.1750 1.3800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        RECT  1.2300 1.1100 1.3500 1.4350 ;
        RECT  0.9300 1.1750 1.3800 1.2950 ;
        RECT  0.8100 1.1700 1.0500 1.2900 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.4740  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5700 1.4300 8.6900 2.2100 ;
        RECT  6.8900 1.5000 8.6900 1.6200 ;
        RECT  0.5550 0.8700 8.4350 0.9900 ;
        RECT  8.3150 0.4000 8.4350 0.9900 ;
        RECT  7.9000 0.8700 8.0500 1.1450 ;
        RECT  7.7300 1.4300 8.0200 1.6200 ;
        RECT  7.9000 0.8700 8.0200 1.6200 ;
        RECT  7.7300 1.4300 7.8500 2.0100 ;
        RECT  7.4750 0.4000 7.5950 0.9900 ;
        RECT  6.8900 1.4300 7.0100 2.0100 ;
        RECT  6.6350 0.4000 6.7550 0.9900 ;
        RECT  5.7350 0.4000 5.8550 0.9900 ;
        RECT  4.8500 0.4000 4.9700 0.9900 ;
        RECT  4.0100 0.4000 4.1300 0.9900 ;
        RECT  3.1700 0.4000 3.2900 0.9900 ;
        RECT  2.3300 0.4000 2.4500 0.9900 ;
        RECT  1.4300 0.4000 1.5500 0.9900 ;
        RECT  0.5550 0.4000 0.6750 0.9900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.7350 -0.1800 8.8550 0.9150 ;
        RECT  7.8950 -0.1800 8.0150 0.7500 ;
        RECT  7.0550 -0.1800 7.1750 0.7500 ;
        RECT  6.1550 -0.1800 6.2750 0.7500 ;
        RECT  5.3150 -0.1800 5.4350 0.7500 ;
        RECT  4.4300 -0.1800 4.5500 0.7500 ;
        RECT  3.5900 -0.1800 3.7100 0.7500 ;
        RECT  2.7500 -0.1800 2.8700 0.7500 ;
        RECT  1.8500 -0.1800 1.9700 0.7500 ;
        RECT  1.0100 -0.1800 1.1300 0.7500 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  1.8500 1.7950 1.9700 2.7900 ;
        RECT  1.0100 1.7950 1.1300 2.7900 ;
        RECT  0.1700 1.4300 0.2900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2700 2.2500 6.4700 2.2500 6.4700 1.6750 5.7500 1.6750 5.7500 2.0100 5.6300 2.0100
                 5.6300 1.6750 4.9100 1.6750 4.9100 2.0100 4.7900 2.0100 4.7900 1.4300 4.9100 1.4300
                 4.9100 1.5550 5.6300 1.5550 5.6300 1.4300 5.7500 1.4300 5.7500 1.5550 6.4700 1.5550
                 6.4700 1.4300 6.5900 1.4300 6.5900 2.1300 7.3100 2.1300 7.3100 1.7400 7.4300 1.7400
                 7.4300 2.1300 8.1500 2.1300 8.1500 1.7400 8.2700 1.7400 ;
        POLYGON  6.1700 2.2500 4.3700 2.2500 4.3700 1.6200 3.6500 1.6200 3.6500 2.0100 3.5300 2.0100
                 3.5300 1.6200 2.8100 1.6200 2.8100 2.0100 2.6900 2.0100 2.6900 1.5000 3.5300 1.5000
                 3.5300 1.4300 3.6500 1.4300 3.6500 1.5000 4.3700 1.5000 4.3700 1.4300 4.4900 1.4300
                 4.4900 2.1300 5.2100 2.1300 5.2100 1.7950 5.3300 1.7950 5.3300 2.1300 6.0500 2.1300
                 6.0500 1.7950 6.1700 1.7950 ;
        POLYGON  4.0700 2.2500 2.2700 2.2500 2.2700 1.6750 1.5500 1.6750 1.5500 2.2100 1.4300 2.2100
                 1.4300 1.6750 0.7100 1.6750 0.7100 2.2100 0.5900 2.2100 0.5900 1.4300 0.7100 1.4300
                 0.7100 1.5550 2.2700 1.5550 2.2700 1.4300 2.3900 1.4300 2.3900 2.1300 3.1100 2.1300
                 3.1100 1.7400 3.2300 1.7400 3.2300 2.1300 3.9500 2.1300 3.9500 1.7400 4.0700 1.7400 ;
    END
END NOR4X6

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1050 1.2600 6.7750 1.3800 ;
        RECT  6.1050 1.2300 6.3650 1.3800 ;
        RECT  6.2450 1.1400 6.3650 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.5050 1.2600 5.2050 1.3800 ;
        RECT  4.9150 1.2300 5.2050 1.3800 ;
        RECT  4.9150 1.1400 5.0350 1.3800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4550 1.2600 3.3550 1.3800 ;
        RECT  3.2350 1.0000 3.3550 1.3800 ;
        RECT  2.6250 1.2300 2.8850 1.3800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1750 1.6700 1.4350 ;
        RECT  1.5350 1.0000 1.6550 1.4350 ;
        RECT  0.7550 1.2800 1.6700 1.4000 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5168  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9750 0.7600 6.9750 0.8800 ;
        RECT  6.8550 0.5900 6.9750 0.8800 ;
        RECT  6.8250 1.5000 6.9450 2.0100 ;
        RECT  2.1300 1.5000 6.9450 1.6200 ;
        RECT  6.0150 0.5900 6.1350 0.8800 ;
        RECT  5.9850 1.5000 6.1050 2.0100 ;
        RECT  5.1750 0.5900 5.2950 0.8800 ;
        RECT  4.3350 0.5900 4.4550 0.8800 ;
        RECT  3.4950 0.5900 3.6150 0.8800 ;
        RECT  2.6550 0.5900 2.7750 0.8800 ;
        RECT  2.1300 0.7600 2.2500 1.6200 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.8150 0.5900 1.9350 0.8800 ;
        RECT  0.9750 0.5900 1.0950 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  7.2750 -0.1800 7.3950 0.6400 ;
        RECT  6.4350 -0.1800 6.5550 0.6400 ;
        RECT  5.5950 -0.1800 5.7150 0.6400 ;
        RECT  4.7550 -0.1800 4.8750 0.6400 ;
        RECT  3.9150 -0.1800 4.0350 0.6400 ;
        RECT  3.0750 -0.1800 3.1950 0.6400 ;
        RECT  2.2350 -0.1800 2.3550 0.6400 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  1.3350 1.9800 1.5750 2.1500 ;
        RECT  1.3350 1.9800 1.4550 2.7900 ;
        RECT  0.4950 1.9800 0.7350 2.1500 ;
        RECT  0.4950 1.9800 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.3650 2.2500 5.5650 2.2500 5.5650 1.8600 4.8450 1.8600 4.8450 2.0100 4.7250 2.0100
                 4.7250 1.8600 4.0050 1.8600 4.0050 2.0100 3.8850 2.0100 3.8850 1.7400 5.6850 1.7400
                 5.6850 2.1300 6.4050 2.1300 6.4050 1.7400 6.5250 1.7400 6.5250 2.1300 7.2450 2.1300
                 7.2450 1.5600 7.3650 1.5600 ;
        POLYGON  5.3250 2.1500 5.2050 2.1500 5.2050 2.2500 2.2950 2.2500 2.2950 2.1500 2.1750 2.1500
                 2.1750 1.9800 2.4150 1.9800 2.4150 2.1300 3.0150 2.1300 3.0150 1.9800 3.2550 1.9800
                 3.2550 2.1300 4.2450 2.1300 4.2450 1.9800 4.4850 1.9800 4.4850 2.1300 5.0850 2.1300
                 5.0850 1.9800 5.3250 1.9800 ;
        POLYGON  3.6150 2.0100 3.4950 2.0100 3.4950 1.8600 2.7750 1.8600 2.7750 2.0100 2.6550 2.0100
                 2.6550 1.8600 1.9350 1.8600 1.9350 2.2100 1.8150 2.2100 1.8150 1.8600 1.0950 1.8600
                 1.0950 2.2100 0.9750 2.2100 0.9750 1.8600 0.2550 1.8600 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.5600 0.2550 1.5600 0.2550 1.7400 0.9750 1.7400 0.9750 1.5600 1.0950 1.5600
                 1.0950 1.7400 1.8150 1.7400 1.8150 1.5600 1.9350 1.5600 1.9350 1.7400 3.6150 1.7400 ;
    END
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4450 0.9400 1.8150 1.1300 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 0.9400 2.5950 1.0900 ;
        RECT  1.2150 1.2500 2.5150 1.3700 ;
        RECT  2.3950 0.9400 2.5150 1.3700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9700 1.4900 2.8350 1.6100 ;
        RECT  2.7150 1.2200 2.8350 1.6100 ;
        RECT  0.9700 1.2800 1.0950 1.6100 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.8550 1.2800 1.0950 1.4000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0200 1.2200 3.2550 1.4600 ;
        RECT  0.4950 1.7300 3.1400 1.8500 ;
        RECT  3.0200 1.2200 3.1400 1.8500 ;
        RECT  2.9700 1.4650 3.1400 1.8500 ;
        RECT  0.4950 1.2200 0.6150 1.8500 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7584  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8550 1.9700 3.4950 2.0900 ;
        RECT  3.3750 0.7000 3.4950 2.0900 ;
        RECT  3.2600 1.7550 3.4950 2.0900 ;
        RECT  0.6150 0.7000 3.4950 0.8200 ;
        RECT  3.0150 0.6500 3.2550 0.8200 ;
        RECT  2.1750 0.6500 2.4150 0.8200 ;
        RECT  1.8550 1.9700 2.0950 2.1500 ;
        RECT  1.3350 0.6500 1.5750 0.8200 ;
        RECT  0.4950 0.6500 0.7350 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.4350 0.4600 3.6750 0.5800 ;
        RECT  3.4350 -0.1800 3.5550 0.5800 ;
        RECT  2.5950 0.4600 2.8350 0.5800 ;
        RECT  2.5950 -0.1800 2.7150 0.5800 ;
        RECT  1.7550 0.4600 1.9950 0.5800 ;
        RECT  1.7550 -0.1800 1.8750 0.5800 ;
        RECT  0.9150 0.4600 1.1550 0.5800 ;
        RECT  0.9150 -0.1800 1.0350 0.5800 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.1950 2.2100 3.4350 2.7900 ;
        RECT  0.4350 1.9700 0.5550 2.7900 ;
        END
    END VDD
END NOR4X2

MACRO NOR4X1
    CLASS CORE ;
    FOREIGN NOR4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.0900 1.6700 1.5750 ;
        RECT  1.5200 1.0900 1.6700 1.5450 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.3050 1.3800 1.7250 ;
        RECT  1.2300 1.0900 1.3500 1.7250 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 1.0300 1.3300 ;
        RECT  0.9100 1.0900 1.0300 1.3300 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.8650 0.5100 1.3400 ;
        RECT  0.0700 0.8650 0.5100 0.9850 ;
        RECT  0.0700 0.8500 0.2200 1.3000 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4572  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7900 0.8850 1.9600 1.1450 ;
        RECT  1.7900 0.8500 1.9100 2.2050 ;
        RECT  0.6500 0.8500 1.9100 0.9700 ;
        RECT  1.4900 0.6800 1.6100 0.9700 ;
        RECT  0.6500 0.6800 0.7700 0.9700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.9100 -0.1800 2.0300 0.7300 ;
        RECT  1.0700 -0.1800 1.1900 0.7300 ;
        RECT  0.2300 -0.1800 0.3500 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  0.4300 1.5550 0.5500 2.7900 ;
        END
    END VDD
END NOR4X1

MACRO NOR4BXL
    CLASS CORE ;
    FOREIGN NOR4BXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0350 0.5350 1.4350 ;
        RECT  0.4150 1.0250 0.5350 1.4350 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9750 1.0950 1.2150 1.2850 ;
        RECT  0.8850 1.1650 1.1450 1.3800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1750 1.6700 1.4350 ;
        RECT  1.3550 1.1750 1.6700 1.2950 ;
        RECT  1.3550 1.0550 1.4750 1.2950 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.1600 2.3050 1.3800 ;
        RECT  2.1150 1.0250 2.2350 1.4100 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2544  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 0.4850 1.6950 0.6050 ;
        RECT  1.4550 0.4850 1.5750 0.9050 ;
        RECT  0.1200 0.7850 1.5750 0.9050 ;
        RECT  0.6750 0.4250 0.7950 0.9050 ;
        RECT  0.5550 1.5550 0.6750 1.7950 ;
        RECT  0.1200 1.5550 0.6750 1.6750 ;
        RECT  0.1200 0.7850 0.2400 1.6750 ;
        RECT  0.0700 0.8850 0.2400 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.9350 -0.1800 2.0550 0.6650 ;
        RECT  1.0950 -0.1800 1.2150 0.6650 ;
        RECT  0.2550 -0.1800 0.3750 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8350 1.5550 1.9550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.5450 1.6500 2.3750 1.6500 2.3750 1.7700 2.2550 1.7700 2.2550 1.5300 2.4250 1.5300
                 2.4250 0.9050 1.8950 0.9050 1.8950 1.0250 1.7750 1.0250 1.7750 0.7850 2.3550 0.7850
                 2.3550 0.4250 2.4750 0.4250 2.4750 0.6650 2.5450 0.6650 ;
    END
END NOR4BXL

MACRO NOR4BX4
    CLASS CORE ;
    FOREIGN NOR4BX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6450 1.2600 7.5650 1.3800 ;
        RECT  6.6450 1.2300 6.9450 1.3800 ;
        RECT  6.6450 1.0000 6.7650 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2350 1.2600 5.8850 1.3800 ;
        RECT  4.9650 1.2300 5.5650 1.3500 ;
        RECT  4.9650 1.0000 5.0850 1.3500 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2050 1.2300 3.7850 1.3500 ;
        RECT  3.2050 1.2300 3.4650 1.3800 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2750 1.0000 0.3950 1.2400 ;
        RECT  0.0700 1.0000 0.3950 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5168  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6450 1.5000 7.7650 2.0100 ;
        RECT  2.9650 1.5000 7.7650 1.6200 ;
        RECT  1.3450 0.7600 7.3450 0.8800 ;
        RECT  7.2250 0.5900 7.3450 0.8800 ;
        RECT  6.8050 1.5000 6.9250 2.0100 ;
        RECT  6.3850 0.5900 6.5050 0.8800 ;
        RECT  5.5450 0.5900 5.6650 0.8800 ;
        RECT  4.7050 0.5900 4.8250 0.8800 ;
        RECT  3.8650 0.5900 3.9850 0.8800 ;
        RECT  2.9150 1.5200 3.1750 1.6700 ;
        RECT  3.0250 0.5900 3.1450 0.8800 ;
        RECT  2.9650 0.7600 3.0850 1.6700 ;
        RECT  2.1850 0.5900 2.3050 0.8800 ;
        RECT  1.3450 0.5900 1.4650 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.6450 -0.1800 7.7650 0.6400 ;
        RECT  6.8050 -0.1800 6.9250 0.6400 ;
        RECT  5.9650 -0.1800 6.0850 0.6400 ;
        RECT  5.1250 -0.1800 5.2450 0.6400 ;
        RECT  4.2850 -0.1800 4.4050 0.6400 ;
        RECT  3.4450 -0.1800 3.5650 0.6400 ;
        RECT  2.6050 -0.1800 2.7250 0.6400 ;
        RECT  1.7650 -0.1800 1.8850 0.6400 ;
        RECT  0.8650 -0.1800 0.9850 0.5300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  2.1250 2.0300 2.3650 2.1500 ;
        RECT  2.1250 2.0300 2.2450 2.7900 ;
        RECT  1.2850 2.0300 1.5250 2.1500 ;
        RECT  1.2850 2.0300 1.4050 2.7900 ;
        RECT  0.1350 1.3600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.1850 2.2500 6.3850 2.2500 6.3850 1.8600 5.7250 1.8600 5.7250 2.0100 5.4850 2.0100
                 5.4850 1.8600 4.8850 1.8600 4.8850 2.0100 4.6450 2.0100 4.6450 1.7400 6.5050 1.7400
                 6.5050 2.1300 7.2250 2.1300 7.2250 1.7400 7.3450 1.7400 7.3450 2.1300 8.0650 2.1300
                 8.0650 1.5600 8.1850 1.5600 ;
        POLYGON  6.1450 2.1500 6.0250 2.1500 6.0250 2.2500 3.0850 2.2500 3.0850 2.1500 2.9650 2.1500
                 2.9650 2.0300 3.2050 2.0300 3.2050 2.1300 3.8050 2.1300 3.8050 2.0300 4.0450 2.0300
                 4.0450 2.1300 5.0650 2.1300 5.0650 1.9800 5.3050 1.9800 5.3050 2.1300 5.9050 2.1300
                 5.9050 1.9800 6.1450 1.9800 ;
        POLYGON  4.4650 2.0100 4.2250 2.0100 4.2250 1.9100 3.6250 1.9100 3.6250 2.0100 3.3850 2.0100
                 3.3850 1.9100 2.7250 1.9100 2.7250 2.2100 2.6050 2.2100 2.6050 1.9100 1.8850 1.9100
                 1.8850 2.2100 1.7650 2.2100 1.7650 1.9100 1.0450 1.9100 1.0450 2.2100 0.9250 2.2100
                 0.9250 1.7900 1.7650 1.7900 1.7650 1.5600 1.8850 1.5600 1.8850 1.7900 2.6050 1.7900
                 2.6050 1.5600 2.7250 1.5600 2.7250 1.7900 3.3850 1.7900 3.3850 1.7400 3.6250 1.7400
                 3.6250 1.7900 4.2250 1.7900 4.2250 1.7400 4.4650 1.7400 ;
        POLYGON  2.1050 1.3200 0.6750 1.3200 0.6750 1.6400 0.5550 1.6400 0.5550 0.6800 0.6750 0.6800
                 0.6750 1.2000 2.1050 1.2000 ;
    END
END NOR4BX4

MACRO NOR4BX2
    CLASS CORE ;
    FOREIGN NOR4BX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.1750 4.1200 1.3850 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2050 1.2300 3.5250 1.4000 ;
        RECT  3.1950 1.1000 3.3550 1.3800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3850 1.2900 2.8850 1.4100 ;
        RECT  2.6250 1.1800 2.8850 1.4100 ;
        RECT  2.3850 1.0000 2.5050 1.4100 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.3950 1.2950 ;
        RECT  0.2750 1.0550 0.3950 1.2950 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7584  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1950 1.5300 4.3150 2.0100 ;
        RECT  2.1450 1.5300 4.3150 1.6500 ;
        RECT  1.3050 0.7600 3.9450 0.8800 ;
        RECT  3.8250 0.5900 3.9450 0.8800 ;
        RECT  2.9850 0.5900 3.1050 0.8800 ;
        RECT  2.1450 0.5900 2.2650 1.6500 ;
        RECT  2.1000 1.1750 2.2650 1.4350 ;
        RECT  1.3050 0.5900 1.4250 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  4.2450 -0.1800 4.3650 0.6400 ;
        RECT  3.4050 -0.1800 3.5250 0.6400 ;
        RECT  2.5650 -0.1800 2.6850 0.6400 ;
        RECT  1.7250 -0.1800 1.8450 0.6400 ;
        RECT  0.8250 -0.1800 0.9450 0.5300 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  1.2250 2.0100 1.4650 2.1500 ;
        RECT  1.2250 2.0100 1.3450 2.7900 ;
        RECT  0.1350 1.5550 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.7350 2.2500 3.7750 2.2500 3.7750 1.8900 3.0550 1.8900 3.0550 2.0100 2.9350 2.0100
                 2.9350 1.7700 3.8950 1.7700 3.8950 2.1300 4.6150 2.1300 4.6150 1.5600 4.7350 1.5600 ;
        POLYGON  3.5350 2.1500 3.4150 2.1500 3.4150 2.2500 2.1850 2.2500 2.1850 2.1500 2.0650 2.1500
                 2.0650 2.0100 2.3050 2.0100 2.3050 2.1300 3.2950 2.1300 3.2950 2.0100 3.5350 2.0100 ;
        POLYGON  2.6650 2.0100 2.5450 2.0100 2.5450 1.8900 1.8250 1.8900 1.8250 2.2100 1.7050 2.2100
                 1.7050 1.8900 0.9850 1.8900 0.9850 2.2100 0.8650 2.2100 0.8650 1.7700 1.7050 1.7700
                 1.7050 1.5600 1.8250 1.5600 1.8250 1.7700 2.6650 1.7700 ;
        POLYGON  1.2250 1.1900 0.6750 1.1900 0.6750 1.6750 0.5550 1.6750 0.5550 0.6800 0.6750 0.6800
                 0.6750 1.0700 1.2250 1.0700 ;
    END
END NOR4BX2

MACRO NOR4BX1
    CLASS CORE ;
    FOREIGN NOR4BX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0000 0.5100 1.4750 ;
        RECT  0.3600 1.0000 0.5100 1.4500 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1650 1.1450 1.4050 ;
        RECT  0.8150 1.0700 1.0550 1.2850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.2100 1.7250 1.3900 ;
        RECT  1.2650 1.2100 1.7250 1.3550 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0600 2.2500 1.5300 ;
        RECT  2.1000 1.0600 2.2200 1.5600 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4572  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 0.5900 1.5750 0.8500 ;
        RECT  0.1200 0.7600 1.5550 0.8800 ;
        RECT  1.4350 0.7300 1.5750 0.8500 ;
        RECT  0.6150 0.5900 0.7350 0.8800 ;
        RECT  0.3950 1.5950 0.5150 2.2100 ;
        RECT  0.1200 1.5950 0.5150 1.7150 ;
        RECT  0.1200 0.7600 0.2400 1.7150 ;
        RECT  0.0700 0.8850 0.2400 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8750 -0.1800 1.9950 0.6400 ;
        RECT  1.0350 -0.1800 1.1550 0.6400 ;
        RECT  0.1950 -0.1800 0.3150 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8050 1.5600 1.9250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4900 1.8000 2.4050 1.8000 2.4050 1.9200 2.2850 1.9200 2.2850 1.6800 2.3700 1.6800
                 2.3700 0.9400 1.9150 0.9400 1.9150 1.0900 1.6750 1.0900 1.6750 0.9700 1.7950 0.9700
                 1.7950 0.8200 2.3550 0.8200 2.3550 0.5900 2.4750 0.5900 2.4750 0.7100 2.4900 0.7100 ;
    END
END NOR4BX1

MACRO NOR4BBXL
    CLASS CORE ;
    FOREIGN NOR4BBXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.1200 0.5650 1.3800 ;
        RECT  0.3050 1.0400 0.5450 1.3800 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.2300 2.8850 1.4450 ;
        RECT  2.5050 1.3250 2.7450 1.5150 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6150 1.2650 1.7350 1.5500 ;
        RECT  1.5200 1.4300 1.6700 1.7250 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9950 1.2400 1.1150 1.6650 ;
        RECT  0.9400 1.3150 1.0900 1.7250 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2544  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0750 1.1750 2.2500 1.4350 ;
        RECT  2.0950 0.4000 2.2150 0.6400 ;
        RECT  1.0750 1.8450 2.1950 1.9650 ;
        RECT  2.0750 0.5200 2.1950 1.9650 ;
        RECT  1.2550 0.7600 2.1950 0.8800 ;
        RECT  1.2550 0.4000 1.3750 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.5150 -0.1800 2.6350 0.6400 ;
        RECT  1.6750 -0.1800 1.7950 0.6400 ;
        RECT  0.7750 -0.1800 0.8950 0.5300 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3150 1.8400 2.4350 2.7900 ;
        RECT  0.1350 1.5000 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1250 1.9000 2.6750 1.9000 2.6750 1.7800 3.0050 1.7800 3.0050 0.9800 2.3150 0.9800
                 2.3150 0.8600 3.0050 0.8600 3.0050 0.6400 2.9350 0.6400 2.9350 0.4000 3.0550 0.4000
                 3.0550 0.5200 3.1250 0.5200 ;
        POLYGON  1.9550 1.1200 0.8050 1.1200 0.8050 1.6200 0.6750 1.6200 0.6750 1.7400 0.5550 1.7400
                 0.5550 1.5000 0.6850 1.5000 0.6850 0.9200 0.5250 0.9200 0.5250 0.6800 0.6450 0.6800
                 0.6450 0.8000 0.8050 0.8000 0.8050 1.0000 1.9550 1.0000 ;
    END
END NOR4BBXL

MACRO NOR4BBX4
    CLASS CORE ;
    FOREIGN NOR4BBX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0100 0.5100 1.4650 ;
        RECT  0.3750 1.0100 0.4950 1.4950 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0100 0.8350 1.3800 ;
        RECT  0.6500 1.0700 0.8000 1.4350 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2900 1.0250 5.4400 1.4800 ;
        RECT  5.3200 1.0000 5.4400 1.4800 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7400 1.1750 7.0550 1.3500 ;
        RECT  6.9350 1.1100 7.0550 1.3500 ;
        RECT  6.7400 1.1750 6.8900 1.4350 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5168  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0550 1.1900 8.1750 2.0100 ;
        RECT  7.2050 1.1900 8.1750 1.3100 ;
        RECT  1.9850 0.7600 7.9850 0.8800 ;
        RECT  7.8650 0.5900 7.9850 0.8800 ;
        RECT  7.2150 1.1750 7.4700 1.4350 ;
        RECT  7.2150 1.1750 7.3350 2.0100 ;
        RECT  7.2050 0.7100 7.3250 1.4300 ;
        RECT  7.0250 0.7100 7.3250 0.8800 ;
        RECT  7.0250 0.5900 7.1450 0.8800 ;
        RECT  6.1850 0.5900 6.3050 0.8800 ;
        RECT  5.3450 0.5900 5.4650 0.8800 ;
        RECT  4.5050 0.5900 4.6250 0.8800 ;
        RECT  3.6650 0.5900 3.7850 0.8800 ;
        RECT  2.8250 0.5900 2.9450 0.8800 ;
        RECT  1.9850 0.5900 2.1050 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.2850 -0.1800 8.4050 0.6400 ;
        RECT  7.4450 -0.1800 7.5650 0.6400 ;
        RECT  6.6050 -0.1800 6.7250 0.6400 ;
        RECT  5.7650 -0.1800 5.8850 0.6400 ;
        RECT  4.9250 -0.1800 5.0450 0.6400 ;
        RECT  4.0850 -0.1800 4.2050 0.6400 ;
        RECT  3.2450 -0.1800 3.3650 0.6400 ;
        RECT  2.4050 -0.1800 2.5250 0.6400 ;
        RECT  1.5650 -0.1800 1.6850 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  2.6250 1.5600 2.7450 2.7900 ;
        RECT  1.7850 1.7200 1.9050 2.7900 ;
        RECT  0.5550 1.6150 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.5950 2.1300 8.5500 2.1300 8.5500 2.2500 5.1150 2.2500 5.1150 1.8400 5.2350 1.8400
                 5.2350 2.1300 5.9550 2.1300 5.9550 1.8400 6.0750 1.8400 6.0750 2.1300 6.7950 2.1300
                 6.7950 1.5550 6.9150 1.5550 6.9150 2.1300 7.6350 2.1300 7.6350 1.4300 7.7550 1.4300
                 7.7550 2.1300 8.4300 2.1300 8.4300 2.0100 8.4750 2.0100 8.4750 1.4300 8.5950 1.4300 ;
        POLYGON  6.4950 2.0100 6.3750 2.0100 6.3750 1.7200 5.6550 1.7200 5.6550 2.0100 5.5350 2.0100
                 5.5350 1.7200 4.4250 1.7200 4.4250 2.0100 4.3050 2.0100 4.3050 1.7200 3.5850 1.7200
                 3.5850 2.0100 3.4650 2.0100 3.4650 1.5600 3.5850 1.5600 3.5850 1.6000 4.3050 1.6000
                 4.3050 1.5600 4.4250 1.5600 4.4250 1.6000 6.3750 1.6000 6.3750 1.4300 6.4950 1.4300 ;
        POLYGON  4.8450 2.2100 4.8000 2.2100 4.8000 2.2500 3.0900 2.2500 3.0900 2.2100 3.0450 2.2100
                 3.0450 1.4400 2.3700 1.4400 2.3700 1.6000 2.3250 1.6000 2.3250 2.2100 2.2050 2.2100
                 2.2050 1.6000 1.4850 1.6000 1.4850 2.2100 1.3650 2.2100 1.3650 1.4800 2.2500 1.4800
                 2.2500 1.3200 3.1650 1.3200 3.1650 2.0900 3.2100 2.0900 3.2100 2.1300 3.8850 2.1300
                 3.8850 1.8400 4.0050 1.8400 4.0050 2.1300 4.6800 2.1300 4.6800 2.0900 4.7250 2.0900
                 4.7250 1.8400 4.8450 1.8400 ;
        POLYGON  3.5850 1.1200 1.7450 1.1200 1.7450 0.8800 1.3250 0.8800 1.3250 0.4800 0.9150 0.4800
                 0.9150 0.8900 0.2400 0.8900 0.2400 1.5850 0.2550 1.5850 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.7050 0.1200 1.7050 0.1200 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000
                 0.2550 0.7700 0.7950 0.7700 0.7950 0.3600 1.4450 0.3600 1.4450 0.7600 1.8650 0.7600
                 1.8650 1.0000 3.5850 1.0000 ;
        POLYGON  1.9050 1.3600 1.1550 1.3600 1.1550 1.4800 1.0950 1.4800 1.0950 2.2100 0.9750 2.2100
                 0.9750 1.3600 1.0350 1.3600 1.0350 0.6000 1.1550 0.6000 1.1550 1.2400 1.9050 1.2400 ;
    END
END NOR4BBX4

MACRO NOR4BBX2
    CLASS CORE ;
    FOREIGN NOR4BBX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 0.9400 0.8550 1.1050 ;
        RECT  0.4950 0.9850 0.6150 1.2650 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 1.3400 1.0950 1.4600 ;
        RECT  0.9750 1.2200 1.0950 1.4600 ;
        RECT  0.5950 1.5200 0.8550 1.6700 ;
        RECT  0.7350 1.3400 0.8550 1.6700 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 1.0450 3.8350 1.4350 ;
        RECT  3.7150 1.0350 3.8350 1.4350 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0750 1.2250 4.7350 1.3500 ;
        RECT  4.0750 1.2250 4.4400 1.3800 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7584  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8550 0.8850 5.1500 1.1450 ;
        RECT  4.8550 0.7100 4.9750 1.6200 ;
        RECT  4.8350 1.5000 4.9550 2.0100 ;
        RECT  2.9950 0.7600 4.9750 0.8800 ;
        RECT  4.6300 0.7100 4.9750 0.8800 ;
        RECT  4.6750 0.5900 4.7950 0.8800 ;
        RECT  3.8350 0.5900 3.9550 0.8800 ;
        RECT  2.0950 0.7000 3.1150 0.7700 ;
        RECT  2.9950 0.5900 3.1150 0.8800 ;
        RECT  2.2150 0.7600 4.9750 0.8200 ;
        RECT  2.0950 0.6500 2.3350 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  5.0950 -0.1800 5.2150 0.6400 ;
        RECT  4.2550 -0.1800 4.3750 0.6400 ;
        RECT  3.4150 -0.1800 3.5350 0.6400 ;
        RECT  2.5150 0.4600 2.7550 0.5800 ;
        RECT  2.5150 -0.1800 2.6350 0.5800 ;
        RECT  1.7350 -0.1800 1.8550 0.6400 ;
        RECT  0.7150 -0.1800 0.8350 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  1.9250 1.6600 2.0450 2.7900 ;
        RECT  0.7150 1.7900 0.8350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.3750 2.1500 5.3300 2.1500 5.3300 2.2500 3.5750 2.2500 3.5750 1.7950 3.6950 1.7950
                 3.6950 2.1300 4.4150 2.1300 4.4150 1.5000 4.5350 1.5000 4.5350 2.1300 5.2100 2.1300
                 5.2100 2.0300 5.2550 2.0300 5.2550 1.5000 5.3750 1.5000 ;
        POLYGON  4.1150 2.0100 3.9950 2.0100 3.9950 1.6750 2.8850 1.6750 2.8850 2.0100 2.7650 2.0100
                 2.7650 1.5550 3.9950 1.5550 3.9950 1.5000 4.1150 1.5000 ;
        POLYGON  3.3050 2.2100 3.2600 2.2100 3.2600 2.2500 2.3450 2.2500 2.3450 1.5400 1.6700 1.5400
                 1.6700 2.0900 1.6250 2.0900 1.6250 2.2100 1.5050 2.2100 1.5050 1.9700 1.5500 1.9700
                 1.5500 1.4200 2.4650 1.4200 2.4650 2.1300 3.1400 2.1300 3.1400 2.0900 3.1850 2.0900
                 3.1850 1.7950 3.3050 1.7950 ;
        POLYGON  2.9150 1.1200 2.6750 1.1200 2.6750 1.0600 1.8550 1.0600 1.8550 0.8800 1.4950 0.8800
                 1.4950 0.4800 1.0750 0.4800 1.0750 0.8200 0.3550 0.8200 0.3550 1.8200 0.2350 1.8200
                 0.2350 0.6000 0.3550 0.6000 0.3550 0.7000 0.9550 0.7000 0.9550 0.3600 1.6150 0.3600
                 1.6150 0.7600 1.9750 0.7600 1.9750 0.9400 2.7950 0.9400 2.7950 1.0000 2.9150 1.0000 ;
        POLYGON  2.0750 1.3000 1.3350 1.3000 1.3350 1.7000 1.3150 1.7000 1.3150 1.8200 1.1950 1.8200
                 1.1950 1.5800 1.2150 1.5800 1.2150 0.8400 1.1950 0.8400 1.1950 0.6000 1.3150 0.6000
                 1.3150 0.7200 1.3350 0.7200 1.3350 1.1800 2.0750 1.1800 ;
    END
END NOR4BBX2

MACRO NOR4BBX1
    CLASS CORE ;
    FOREIGN NOR4BBX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2450 1.0200 0.3650 1.2600 ;
        RECT  0.0700 1.0200 0.3650 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.2500 2.8900 1.5000 ;
        RECT  2.6250 1.2300 2.8850 1.5000 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.5200 1.3400 1.6400 1.7250 ;
        RECT  1.4300 1.2200 1.5500 1.4600 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9950 1.2200 1.1150 1.4600 ;
        RECT  0.9400 1.4650 1.0900 1.7250 ;
        RECT  0.9700 1.3400 1.0900 1.7250 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4572  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0700 1.4650 2.2500 1.7250 ;
        RECT  1.3150 0.7100 2.2150 0.8300 ;
        RECT  2.0950 0.5900 2.2150 0.8300 ;
        RECT  0.9500 1.8450 2.1900 1.9650 ;
        RECT  2.0700 0.7100 2.1900 1.9650 ;
        RECT  1.1950 0.6500 1.4350 0.7700 ;
        RECT  0.9500 1.8450 1.0700 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.5150 -0.1800 2.6350 0.8300 ;
        RECT  1.6150 0.4600 1.8550 0.5800 ;
        RECT  1.6150 -0.1800 1.7350 0.5800 ;
        RECT  0.7750 -0.1800 0.8950 0.5300 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3100 1.8450 2.4300 2.7900 ;
        RECT  0.1350 1.9800 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1300 1.7400 2.9700 1.7400 2.9700 1.8600 2.8500 1.8600 2.8500 1.6200 3.0100 1.6200
                 3.0100 1.1100 2.3100 1.1100 2.3100 0.9900 2.9350 0.9900 2.9350 0.5900 3.0550 0.5900
                 3.0550 0.8700 3.1300 0.8700 ;
        POLYGON  1.9500 1.1000 0.6800 1.1000 0.6800 1.5800 0.5600 1.5800 0.5600 0.9800 0.5250 0.9800
                 0.5250 0.6800 0.6450 0.6800 0.6450 0.8600 0.6800 0.8600 0.6800 0.9800 1.9500 0.9800 ;
    END
END NOR4BBX1

MACRO NOR3XL
    CLASS CORE ;
    FOREIGN NOR3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 1.2800 0.8200 1.7550 ;
        RECT  0.6500 1.2800 0.8200 1.7300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3500 1.3400 0.5300 1.7250 ;
        RECT  0.3600 1.3300 0.5100 1.7250 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0500 1.2800 1.1700 1.6500 ;
        RECT  0.9400 1.3600 1.0900 1.7250 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2448  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5700 1.0400 1.5300 1.1600 ;
        RECT  1.4100 0.6800 1.5300 1.1600 ;
        RECT  1.2900 0.8850 1.4100 1.8900 ;
        RECT  1.2100 1.7700 1.3300 2.0100 ;
        RECT  1.2300 0.8850 1.5300 1.1600 ;
        RECT  0.5700 0.6800 0.6900 1.1600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9900 -0.1800 1.1100 0.9200 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.2200 1.8450 0.3400 2.7900 ;
        END
    END VDD
END NOR3XL

MACRO NOR3X8
    CLASS CORE ;
    FOREIGN NOR3X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6950 0.8100 9.8150 1.2100 ;
        RECT  9.0050 0.8100 9.8150 0.9300 ;
        RECT  1.8550 0.7300 9.1250 0.8450 ;
        RECT  6.0350 0.8100 9.8150 0.8500 ;
        RECT  7.1500 1.0300 7.3900 1.1500 ;
        RECT  7.1500 0.7300 7.2700 1.1500 ;
        RECT  1.8550 0.7250 6.1550 0.8450 ;
        RECT  4.4650 1.0300 4.7050 1.1500 ;
        RECT  4.5850 0.7250 4.7050 1.1500 ;
        RECT  1.8550 0.7250 2.0150 1.0900 ;
        RECT  1.7350 1.0350 1.9750 1.1550 ;
        RECT  1.7550 0.9400 2.0150 1.0900 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 1.2300 9.5550 1.3800 ;
        RECT  9.2950 1.0500 9.5350 1.3800 ;
        RECT  8.7650 1.0500 9.5350 1.1700 ;
        RECT  7.9700 0.9700 8.8850 1.0900 ;
        RECT  7.6500 1.0500 8.1550 1.1700 ;
        RECT  6.8550 1.2700 7.7700 1.3900 ;
        RECT  7.6500 1.0500 7.7700 1.3900 ;
        RECT  6.8550 1.0500 6.9750 1.3900 ;
        RECT  5.7950 1.0500 6.9750 1.1700 ;
        RECT  5.1950 0.9650 5.9150 1.0850 ;
        RECT  4.8250 1.0500 5.3150 1.1700 ;
        RECT  4.2250 1.2700 4.9450 1.3900 ;
        RECT  4.8250 1.0500 4.9450 1.3900 ;
        RECT  4.2250 0.9900 4.3450 1.3900 ;
        RECT  3.6950 0.9900 4.3450 1.1100 ;
        RECT  3.6950 0.9650 3.8150 1.2300 ;
        RECT  2.9000 0.9650 3.8150 1.0850 ;
        RECT  2.1350 1.0550 3.0200 1.1750 ;
        RECT  1.4050 1.2750 2.2550 1.3950 ;
        RECT  2.1350 1.0550 2.2550 1.3950 ;
        RECT  1.4050 1.0550 1.5250 1.3950 ;
        RECT  0.7550 1.0550 1.5250 1.1750 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.3150 1.2100 8.5550 1.3300 ;
        RECT  8.3150 1.2100 8.4350 1.6300 ;
        RECT  2.5650 1.5100 8.4350 1.6300 ;
        RECT  5.4350 1.2050 5.6750 1.3250 ;
        RECT  5.4350 1.2050 5.5550 1.6300 ;
        RECT  3.3550 1.2050 3.4750 1.6300 ;
        RECT  3.2350 1.2050 3.4750 1.3250 ;
        RECT  0.9750 1.5150 2.6850 1.6350 ;
        RECT  0.9750 1.2950 1.0950 1.6350 ;
        RECT  0.4450 1.2950 1.0950 1.4150 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        RECT  0.4450 1.1250 0.5650 1.4150 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.6308  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4950 0.4850 10.3350 0.6050 ;
        RECT  9.8350 1.5200 10.1350 1.6700 ;
        RECT  1.8350 1.7550 10.0550 1.8750 ;
        RECT  9.9350 0.4850 10.0550 1.8750 ;
        RECT  9.8350 1.4700 9.9550 2.2100 ;
        RECT  7.4900 1.7500 7.6100 2.2100 ;
        RECT  4.2450 1.7500 4.3650 2.2100 ;
        RECT  1.8350 1.7550 1.9550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  9.6150 -0.1800 9.8550 0.3650 ;
        RECT  8.6550 -0.1800 8.8950 0.3650 ;
        RECT  7.6950 -0.1800 7.9350 0.3650 ;
        RECT  6.7350 -0.1800 6.9750 0.3650 ;
        RECT  5.7750 -0.1800 6.0150 0.3650 ;
        RECT  4.8150 -0.1800 5.0550 0.3650 ;
        RECT  3.8550 -0.1800 4.0950 0.3650 ;
        RECT  2.8950 -0.1800 3.1350 0.3650 ;
        RECT  1.9350 -0.1800 2.1750 0.3650 ;
        RECT  0.9750 -0.1800 1.2150 0.3650 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  8.5950 1.9950 8.8350 2.1500 ;
        RECT  8.5950 1.9950 8.7150 2.7900 ;
        RECT  5.5150 1.9950 5.7550 2.1500 ;
        RECT  5.5150 1.9950 5.6350 2.7900 ;
        RECT  2.9550 1.9950 3.1950 2.1500 ;
        RECT  2.9550 1.9950 3.0750 2.7900 ;
        RECT  0.3350 1.5350 0.4550 2.7900 ;
        END
    END VDD
END NOR3X8

MACRO NOR3X6
    CLASS CORE ;
    FOREIGN NOR3X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9050 1.0550 7.1450 1.1750 ;
        RECT  6.9050 0.8200 7.0250 1.1750 ;
        RECT  4.7850 0.8200 7.0250 0.9400 ;
        RECT  3.9800 1.0350 4.9050 1.1550 ;
        RECT  4.7850 0.8200 4.9050 1.1550 ;
        RECT  4.2450 1.0350 4.4850 1.1750 ;
        RECT  3.9800 0.8200 4.1000 1.1550 ;
        RECT  2.3900 0.8200 4.1000 0.9400 ;
        RECT  2.3900 0.8200 2.5100 1.0900 ;
        RECT  1.7550 0.9700 2.5100 1.0900 ;
        RECT  1.7550 0.9400 2.0150 1.0900 ;
        RECT  1.7400 1.0550 1.9800 1.1750 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.2300 7.5250 1.3800 ;
        RECT  6.5250 1.2950 7.4800 1.4150 ;
        RECT  7.3600 1.0200 7.4800 1.4150 ;
        RECT  5.9950 1.2800 6.6600 1.4000 ;
        RECT  5.9950 1.0600 6.1150 1.4000 ;
        RECT  5.2000 1.0600 6.1150 1.1800 ;
        RECT  5.2000 1.0600 5.3200 1.4150 ;
        RECT  4.7500 1.2750 5.3200 1.3950 ;
        RECT  3.4250 1.2950 4.8700 1.4150 ;
        RECT  3.6900 1.1750 3.8100 1.4150 ;
        RECT  3.4250 1.0600 3.5450 1.4150 ;
        RECT  2.6300 1.0600 3.5450 1.1800 ;
        RECT  2.6300 1.0600 2.7500 1.4000 ;
        RECT  2.1000 1.2800 2.7500 1.4000 ;
        RECT  1.3050 1.2950 2.2200 1.4150 ;
        RECT  1.3050 1.0800 1.4250 1.4150 ;
        RECT  0.7550 1.0800 1.4250 1.2000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7000 1.1050 7.8200 1.3450 ;
        RECT  7.7000 1.1050 7.7650 1.6200 ;
        RECT  0.9750 1.5350 7.7200 1.6550 ;
        RECT  7.6000 1.5000 7.7650 1.6200 ;
        RECT  7.6450 1.2250 7.7200 1.6550 ;
        RECT  5.4800 1.3000 5.7200 1.6550 ;
        RECT  2.9750 1.3000 3.2150 1.6550 ;
        RECT  0.9750 1.3200 1.0950 1.6550 ;
        RECT  0.4450 1.3200 1.0950 1.4400 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        RECT  0.4450 1.2000 0.5650 1.4400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.9271  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8400 1.7750 8.0600 1.8950 ;
        RECT  7.9400 0.5800 8.0600 1.8950 ;
        RECT  7.9000 1.4650 8.0600 1.8950 ;
        RECT  0.5550 0.5800 8.0600 0.7000 ;
        RECT  7.2800 0.4000 7.4000 0.9000 ;
        RECT  6.9600 1.7750 7.0800 2.2100 ;
        RECT  6.3200 0.4000 6.4400 0.7000 ;
        RECT  5.3600 0.4000 5.4800 0.7000 ;
        RECT  4.5850 1.7750 4.7050 2.2100 ;
        RECT  4.4000 0.4000 4.5200 0.9150 ;
        RECT  3.4400 0.4000 3.5600 0.7000 ;
        RECT  2.4800 0.4000 2.6000 0.7000 ;
        RECT  1.8400 1.7750 1.9600 2.2100 ;
        RECT  1.5150 0.4000 1.6350 0.9150 ;
        RECT  0.5550 0.4000 0.6750 0.9200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  6.7400 0.3400 6.9800 0.4600 ;
        RECT  6.7400 -0.1800 6.8600 0.4600 ;
        RECT  5.7800 0.3400 6.0200 0.4600 ;
        RECT  5.7800 -0.1800 5.9000 0.4600 ;
        RECT  4.8200 0.3400 5.0600 0.4600 ;
        RECT  4.8200 -0.1800 4.9400 0.4600 ;
        RECT  3.8600 0.3400 4.1000 0.4600 ;
        RECT  3.8600 -0.1800 3.9800 0.4600 ;
        RECT  2.9000 0.3400 3.1400 0.4600 ;
        RECT  2.9000 -0.1800 3.0200 0.4600 ;
        RECT  1.9400 0.3400 2.1800 0.4600 ;
        RECT  1.9400 -0.1800 2.0600 0.4600 ;
        RECT  0.9750 0.3400 1.2150 0.4600 ;
        RECT  0.9750 -0.1800 1.0950 0.4600 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.8000 2.0150 8.0400 2.1500 ;
        RECT  7.8000 2.0150 7.9200 2.7900 ;
        RECT  5.7600 2.0150 6.0000 2.1500 ;
        RECT  5.7600 2.0150 5.8800 2.7900 ;
        RECT  2.7400 2.0150 2.9800 2.1500 ;
        RECT  2.7400 2.0150 2.8600 2.7900 ;
        RECT  0.3350 1.5600 0.4550 2.7900 ;
        END
    END VDD
END NOR3X6

MACRO NOR3X4
    CLASS CORE ;
    FOREIGN NOR3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0550 0.9700 4.2950 1.0900 ;
        RECT  4.0550 0.8200 4.1750 1.0900 ;
        RECT  1.8550 0.8200 4.1750 0.9400 ;
        RECT  1.7350 0.9700 2.0150 1.0900 ;
        RECT  1.7550 0.9400 2.0150 1.0900 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8750 1.0100 4.9950 1.2500 ;
        RECT  4.7100 1.0100 4.9950 1.1450 ;
        RECT  4.7100 0.8850 4.8600 1.1450 ;
        RECT  3.5950 1.2100 4.7300 1.3300 ;
        RECT  4.6100 1.0250 4.7300 1.3300 ;
        RECT  3.5950 1.0600 3.7150 1.3300 ;
        RECT  2.8000 1.0600 3.7150 1.1800 ;
        RECT  2.2550 1.0700 2.9200 1.1900 ;
        RECT  1.4750 1.2100 2.3900 1.3300 ;
        RECT  2.2550 1.0700 2.3900 1.3300 ;
        RECT  1.4750 1.0800 1.5950 1.3300 ;
        RECT  0.9750 1.0800 1.5950 1.2000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9200 1.4500 5.3350 1.5700 ;
        RECT  5.2150 1.2400 5.3350 1.5700 ;
        RECT  3.0950 1.3000 3.3350 1.5700 ;
        RECT  0.9200 1.3200 1.0400 1.5700 ;
        RECT  0.3900 1.3200 1.0400 1.4400 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2416  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.4550 1.4650 5.7300 1.7250 ;
        RECT  1.8350 1.6900 5.5750 1.8100 ;
        RECT  5.4550 0.5800 5.5750 1.8100 ;
        RECT  0.4950 0.5800 5.5750 0.7000 ;
        RECT  4.3950 1.6900 4.5150 2.2100 ;
        RECT  1.8350 1.6900 1.9550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.7750 0.3400 6.0150 0.4600 ;
        RECT  5.7750 -0.1800 5.8950 0.4600 ;
        RECT  4.8150 0.3400 5.0550 0.4600 ;
        RECT  4.8150 -0.1800 4.9350 0.4600 ;
        RECT  3.8550 0.3400 4.0950 0.4600 ;
        RECT  3.8550 -0.1800 3.9750 0.4600 ;
        RECT  2.8950 0.3400 3.1350 0.4600 ;
        RECT  2.8950 -0.1800 3.0150 0.4600 ;
        RECT  1.9350 0.3400 2.1750 0.4600 ;
        RECT  1.9350 -0.1800 2.0550 0.4600 ;
        RECT  0.9750 0.3400 1.2150 0.4600 ;
        RECT  0.9750 -0.1800 1.0950 0.4600 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.2950 1.9300 5.5350 2.1500 ;
        RECT  5.2950 1.9300 5.4150 2.7900 ;
        RECT  2.9550 1.9300 3.1950 2.1500 ;
        RECT  2.9550 1.9300 3.0750 2.7900 ;
        RECT  0.5550 1.5600 0.6750 2.7900 ;
        END
    END VDD
END NOR3X4

MACRO NOR3X2
    CLASS CORE ;
    FOREIGN NOR3X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5550 0.8200 2.6750 1.1500 ;
        RECT  0.3900 0.8200 2.6750 0.9400 ;
        RECT  0.3900 0.8200 0.5100 1.1500 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0600 2.3350 1.3000 ;
        RECT  2.1000 1.0600 2.2500 1.4350 ;
        RECT  0.9750 1.0600 2.3350 1.1800 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6050 1.3000 1.8450 1.4200 ;
        RECT  1.4650 1.5200 1.7250 1.6700 ;
        RECT  1.6050 1.3000 1.7250 1.6700 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6208  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7950 0.5950 3.1200 0.8550 ;
        RECT  1.7350 1.7900 2.9150 1.9100 ;
        RECT  2.7950 0.5800 2.9150 1.9100 ;
        RECT  0.4950 0.5800 2.9150 0.7000 ;
        RECT  1.7350 1.7900 1.8550 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.8950 0.3400 3.1350 0.4600 ;
        RECT  2.8950 -0.1800 3.0150 0.4600 ;
        RECT  1.9350 0.3400 2.1750 0.4600 ;
        RECT  1.9350 -0.1800 2.0550 0.4600 ;
        RECT  0.9750 0.3400 1.2150 0.4600 ;
        RECT  0.9750 -0.1800 1.0950 0.4600 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.6350 2.0300 2.8750 2.1500 ;
        RECT  2.6350 2.0300 2.7550 2.7900 ;
        RECT  0.5550 1.5600 0.6750 2.7900 ;
        END
    END VDD
END NOR3X2

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0000 0.8000 1.4550 ;
        RECT  0.6500 1.0000 0.7700 1.4800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.8850 0.5100 1.2900 ;
        RECT  0.3300 0.9100 0.4500 1.3300 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 1.1300 1.1100 1.5550 ;
        RECT  0.9400 1.1750 1.0900 1.5800 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 0.7600 1.5150 0.8800 ;
        RECT  1.3950 0.5900 1.5150 0.8800 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        RECT  1.2300 0.7600 1.3500 2.1000 ;
        RECT  0.5550 0.6450 0.8550 0.7650 ;
        RECT  0.5550 0.5250 0.6750 0.7650 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.1700 1.4500 0.2900 2.7900 ;
        END
    END VDD
END NOR3X1

MACRO NOR3BXL
    CLASS CORE ;
    FOREIGN NOR3BXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0000 0.5100 1.5000 ;
        RECT  0.3600 1.0000 0.5100 1.4700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.9350 1.4000 ;
        RECT  0.8150 1.1600 0.9350 1.4000 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.1500 1.7250 1.3800 ;
        RECT  1.4750 1.0900 1.5950 1.5000 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2448  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9150 0.4600 1.1550 0.5800 ;
        RECT  0.1200 0.7600 1.0350 0.8800 ;
        RECT  0.9150 0.4600 1.0350 0.8800 ;
        RECT  0.3350 1.6200 0.4550 1.8600 ;
        RECT  0.1200 1.6200 0.4550 1.7400 ;
        RECT  0.1350 0.4000 0.2550 0.8800 ;
        RECT  0.1200 0.7600 0.2400 1.7400 ;
        RECT  0.0700 0.8850 0.2400 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.2950 1.6200 1.4150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9650 1.6200 1.8350 1.6200 1.8350 1.7400 1.7150 1.7400 1.7150 1.5000 1.8450 1.5000
                 1.8450 0.9700 1.3450 0.9700 1.3450 1.0600 1.2250 1.0600 1.2250 0.8200 1.3450 0.8200
                 1.3450 0.8500 1.8450 0.8500 1.8450 0.6400 1.8150 0.6400 1.8150 0.4000 1.9350 0.4000
                 1.9350 0.5200 1.9650 0.5200 ;
    END
END NOR3BXL

MACRO NOR3BX4
    CLASS CORE ;
    FOREIGN NOR3BX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1800 0.9700 4.4200 1.0900 ;
        RECT  4.1800 0.8200 4.3000 1.0900 ;
        RECT  2.8400 0.8200 4.3000 0.9400 ;
        RECT  1.8600 0.9700 2.9600 1.0900 ;
        RECT  2.8400 0.8200 2.9600 1.0900 ;
        RECT  2.0450 0.9400 2.3050 1.0900 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9200 0.9900 6.1600 1.2000 ;
        RECT  5.8150 0.9300 6.0750 1.1600 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6300 1.0800 5.4000 1.2000 ;
        RECT  3.7200 1.2100 4.7500 1.3300 ;
        RECT  4.6300 1.0800 4.7500 1.3300 ;
        RECT  3.7200 1.0600 3.8400 1.3300 ;
        RECT  3.0800 1.0600 3.8400 1.1800 ;
        RECT  0.9400 1.2100 3.2000 1.3300 ;
        RECT  3.0800 1.0600 3.2000 1.3300 ;
        RECT  0.9400 0.8850 1.0900 1.3300 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2416  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.5800 5.6600 0.7000 ;
        RECT  4.2000 1.6900 4.3200 2.2100 ;
        RECT  0.3600 1.6900 4.3200 1.8100 ;
        RECT  1.6400 1.6900 1.7600 2.2100 ;
        RECT  0.3600 0.5800 0.4800 1.8100 ;
        RECT  0.0700 1.4650 0.4800 1.5850 ;
        RECT  0.0700 1.4650 0.2200 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  5.9000 -0.1800 6.0200 0.6400 ;
        RECT  4.9400 0.3400 5.1800 0.4600 ;
        RECT  4.9400 -0.1800 5.0600 0.4600 ;
        RECT  3.9800 0.3400 4.2200 0.4600 ;
        RECT  3.9800 -0.1800 4.1000 0.4600 ;
        RECT  3.0200 0.3400 3.2600 0.4600 ;
        RECT  3.0200 -0.1800 3.1400 0.4600 ;
        RECT  2.0600 0.3400 2.3000 0.4600 ;
        RECT  2.0600 -0.1800 2.1800 0.4600 ;
        RECT  1.1000 0.3400 1.3400 0.4600 ;
        RECT  1.1000 -0.1800 1.2200 0.4600 ;
        RECT  0.1400 0.3400 0.3800 0.4600 ;
        RECT  0.1400 -0.1800 0.2600 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  5.7000 1.5600 5.8200 2.7900 ;
        RECT  3.0400 1.9300 3.2800 2.1500 ;
        RECT  3.0400 1.9300 3.1600 2.7900 ;
        RECT  0.4000 1.9300 0.6400 2.1500 ;
        RECT  0.4000 1.9300 0.5200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.5000 0.7700 6.4000 0.7700 6.4000 1.5600 6.2400 1.5600 6.2400 2.2100 6.1200 2.2100
                 6.1200 1.4400 5.4150 1.4400 5.4150 1.5700 0.6000 1.5700 0.6000 1.2400 0.7200 1.2400
                 0.7200 1.4500 3.3200 1.4500 3.3200 1.3000 3.5600 1.3000 3.5600 1.4500 5.2950 1.4500
                 5.2950 1.3200 5.5200 1.3200 5.5200 1.2800 5.7600 1.2800 5.7600 1.3200 6.2800 1.3200
                 6.2800 0.7700 6.2600 0.7700 6.2600 0.6500 6.5000 0.6500 ;
    END
END NOR3BX4

MACRO NOR3BX2
    CLASS CORE ;
    FOREIGN NOR3BX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.8850 1.1750 3.1600 1.4150 ;
        RECT  2.8850 1.1750 3.1200 1.4350 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0600 2.4000 1.3000 ;
        RECT  2.1000 1.0600 2.2500 1.4350 ;
        RECT  0.8200 1.0600 2.4000 1.1800 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.8100 1.3000 1.9300 1.7250 ;
        RECT  1.6900 1.3000 1.9300 1.4200 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6338  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3000 0.5800 2.7200 0.7000 ;
        RECT  1.4500 1.3000 1.5700 2.2100 ;
        RECT  0.0700 1.3000 1.5700 1.4200 ;
        RECT  0.0700 1.1750 0.4200 1.4200 ;
        RECT  0.3000 0.5800 0.4200 1.4200 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  2.9600 -0.1800 3.0800 0.7000 ;
        RECT  2.0000 0.3400 2.2400 0.4600 ;
        RECT  2.0000 -0.1800 2.1200 0.4600 ;
        RECT  1.0400 0.3400 1.2800 0.4600 ;
        RECT  1.0400 -0.1800 1.1600 0.4600 ;
        RECT  0.0800 0.3400 0.3200 0.4600 ;
        RECT  0.0800 -0.1800 0.2000 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  2.7600 1.5600 2.8800 2.7900 ;
        RECT  0.4000 1.5600 0.5200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.5000 0.7000 3.4000 0.7000 3.4000 1.6550 3.3600 1.6550 3.3600 1.8000 3.2400 1.8000
                 3.2400 1.5350 3.2800 1.5350 3.2800 0.9400 2.7200 0.9400 2.7200 1.1700 2.6000 1.1700
                 2.6000 0.9400 0.6600 0.9400 0.6600 1.1500 0.5400 1.1500 0.5400 0.8200 3.2800 0.8200
                 3.2800 0.5800 3.3800 0.5800 3.3800 0.4600 3.5000 0.4600 ;
    END
END NOR3BX2

MACRO NOR3BX1
    CLASS CORE ;
    FOREIGN NOR3BX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0000 0.5100 1.4700 ;
        RECT  0.3600 1.0000 0.4800 1.5000 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9250 1.1650 1.0900 1.4350 ;
        RECT  0.8550 1.0300 0.9900 1.2850 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5750 1.0000 1.6950 1.4900 ;
        RECT  1.5200 1.0000 1.6950 1.4600 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 0.7600 1.0950 0.8800 ;
        RECT  0.9750 0.5900 1.0950 0.8800 ;
        RECT  0.3750 1.6200 0.4950 2.2100 ;
        RECT  0.1200 1.6200 0.4950 1.7400 ;
        RECT  0.1350 0.5900 0.2550 0.8800 ;
        RECT  0.1200 0.7600 0.2400 1.7400 ;
        RECT  0.0700 1.1750 0.2400 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.3350 1.5800 1.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 1.8500 1.8150 1.8500 1.8150 0.8800 1.3550 0.8800 1.3550 1.1700 1.2350 1.1700
                 1.2350 0.7600 1.8150 0.7600 1.8150 0.4000 1.9350 0.4000 ;
    END
END NOR3BX1

MACRO NOR2XL
    CLASS CORE ;
    FOREIGN NOR2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.1600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.0250 0.6750 1.2650 ;
        RECT  0.3900 1.1450 0.6750 1.2650 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 0.7900 0.2400 1.2250 ;
        RECT  0.0700 0.7300 0.2200 1.1450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1776  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7950 0.7850 0.9150 1.8250 ;
        RECT  0.6500 1.4650 0.9150 1.7250 ;
        RECT  0.4950 0.7850 0.9150 0.9050 ;
        RECT  0.4950 0.6650 0.6150 0.9050 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.1600 0.1800 ;
        RECT  0.9050 -0.1800 1.0250 0.3850 ;
        RECT  0.1350 -0.1800 0.2550 0.3850 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.1600 2.7900 ;
        RECT  0.1550 1.7050 0.2750 2.7900 ;
        END
    END VDD
END NOR2XL

MACRO NOR2X8
    CLASS CORE ;
    FOREIGN NOR2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8550 1.0500 5.0950 1.1700 ;
        RECT  0.6800 0.9650 4.9750 1.0850 ;
        RECT  3.4950 0.9650 3.7350 1.1700 ;
        RECT  1.9950 0.9650 2.2350 1.1700 ;
        RECT  0.6500 1.0550 0.8000 1.4350 ;
        RECT  0.4350 1.0550 0.8000 1.1750 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3750 1.1900 5.8350 1.3100 ;
        RECT  1.3150 1.2900 5.4950 1.4100 ;
        RECT  5.2350 1.2300 5.8350 1.3100 ;
        RECT  3.9950 1.2100 4.2350 1.4100 ;
        RECT  2.7350 1.2050 2.9750 1.4100 ;
        RECT  1.1950 1.2050 1.4350 1.3250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0216  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.5300 6.0750 1.6500 ;
        RECT  5.9550 0.7100 6.0750 1.6500 ;
        RECT  5.8150 1.4700 6.0200 1.7250 ;
        RECT  5.8700 1.4650 6.0750 1.6500 ;
        RECT  0.4950 0.7100 6.0750 0.8300 ;
        RECT  5.8150 1.4700 5.9350 2.2100 ;
        RECT  4.3350 1.5300 4.4550 2.2100 ;
        RECT  2.5350 1.5300 2.6550 2.2100 ;
        RECT  1.1750 1.5300 1.2950 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.9550 0.4600 6.1950 0.5800 ;
        RECT  5.9550 -0.1800 6.0750 0.5800 ;
        RECT  5.1150 0.4600 5.3550 0.5800 ;
        RECT  5.1150 -0.1800 5.2350 0.5800 ;
        RECT  4.2750 0.4600 4.5150 0.5800 ;
        RECT  4.2750 -0.1800 4.3950 0.5800 ;
        RECT  3.4350 0.4600 3.6750 0.5800 ;
        RECT  3.4350 -0.1800 3.5550 0.5800 ;
        RECT  2.5950 0.4600 2.8350 0.5800 ;
        RECT  2.5950 -0.1800 2.7150 0.5800 ;
        RECT  1.7550 0.4600 1.9950 0.5800 ;
        RECT  1.7550 -0.1800 1.8750 0.5800 ;
        RECT  0.9150 0.4600 1.1550 0.5800 ;
        RECT  0.9150 -0.1800 1.0350 0.5800 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.1750 1.7700 5.2950 2.7900 ;
        RECT  3.2950 1.7700 3.4150 2.7900 ;
        RECT  1.8950 1.7700 2.0150 2.7900 ;
        RECT  0.3350 1.4650 0.4550 2.7900 ;
        END
    END VDD
END NOR2X8

MACRO NOR2X6
    CLASS CORE ;
    FOREIGN NOR2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4150 0.9900 4.5350 1.2600 ;
        RECT  0.6800 0.9900 4.5350 1.1100 ;
        RECT  3.1750 0.9900 3.4150 1.1950 ;
        RECT  1.9550 0.9900 2.1950 1.1950 ;
        RECT  0.6500 1.0800 0.8000 1.4350 ;
        RECT  0.4350 1.0800 0.8000 1.2000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.3000 4.2350 1.4200 ;
        RECT  3.7850 1.2300 4.0450 1.4200 ;
        RECT  1.3150 1.3150 3.9050 1.4350 ;
        RECT  2.3150 1.3000 2.5550 1.4350 ;
        RECT  1.1950 1.3000 1.4350 1.4200 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.4496  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.5550 4.7750 1.6750 ;
        RECT  4.6550 0.7500 4.7750 1.6750 ;
        RECT  4.4200 1.4650 4.7750 1.6750 ;
        RECT  0.5550 0.7500 4.7750 0.8700 ;
        RECT  4.4200 1.4650 4.5700 1.7250 ;
        RECT  3.9350 1.5550 4.0550 2.2100 ;
        RECT  3.9150 0.4000 4.0350 0.8700 ;
        RECT  3.0750 0.4000 3.1950 0.8700 ;
        RECT  2.4950 1.5550 2.6150 2.2100 ;
        RECT  2.2350 0.4000 2.3550 0.8700 ;
        RECT  1.3950 0.4000 1.5150 0.8700 ;
        RECT  1.1750 1.5550 1.2950 2.2100 ;
        RECT  0.5550 0.4000 0.6750 0.8700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  4.2750 0.4600 4.5150 0.6300 ;
        RECT  4.2750 -0.1800 4.3950 0.6300 ;
        RECT  3.4350 0.4600 3.6750 0.6300 ;
        RECT  3.4350 -0.1800 3.5550 0.6300 ;
        RECT  2.5950 0.4600 2.8350 0.6300 ;
        RECT  2.5950 -0.1800 2.7150 0.6300 ;
        RECT  1.7550 0.4600 1.9950 0.6300 ;
        RECT  1.7550 -0.1800 1.8750 0.6300 ;
        RECT  0.9150 0.4600 1.1550 0.6300 ;
        RECT  0.9150 -0.1800 1.0350 0.6300 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  4.5750 1.8450 4.6950 2.7900 ;
        RECT  3.2950 1.7950 3.4150 2.7900 ;
        RECT  1.8150 1.7950 1.9350 2.7900 ;
        RECT  0.3350 1.5600 0.4550 2.7900 ;
        END
    END VDD
END NOR2X6

MACRO NOR2X4
    CLASS CORE ;
    FOREIGN NOR2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4150 0.9900 3.3350 1.1100 ;
        RECT  1.6950 0.9900 1.9350 1.1300 ;
        RECT  0.6500 0.9900 0.8000 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1950 1.2600 2.5950 1.3800 ;
        RECT  2.3350 1.2300 2.5950 1.3800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9664  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2750 1.5000 3.5750 1.6200 ;
        RECT  3.4550 0.7300 3.5750 1.6200 ;
        RECT  3.2050 1.2300 3.5750 1.3800 ;
        RECT  0.5550 0.7300 3.5750 0.8500 ;
        RECT  3.0750 0.6100 3.1950 0.8500 ;
        RECT  2.5550 1.5000 2.6750 2.2100 ;
        RECT  2.2350 0.6100 2.3550 0.8500 ;
        RECT  1.3950 0.6100 1.5150 0.8500 ;
        RECT  1.2750 1.5000 1.3950 2.2100 ;
        RECT  0.5550 0.6100 0.6750 0.8500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.4350 0.4800 3.6750 0.6000 ;
        RECT  3.4350 -0.1800 3.5550 0.6000 ;
        RECT  2.5950 0.4800 2.8350 0.6000 ;
        RECT  2.5950 -0.1800 2.7150 0.6000 ;
        RECT  1.7550 0.4800 1.9950 0.6000 ;
        RECT  1.7550 -0.1800 1.8750 0.6000 ;
        RECT  0.9150 0.4800 1.1550 0.6000 ;
        RECT  0.9150 -0.1800 1.0350 0.6000 ;
        RECT  0.1350 -0.1800 0.2550 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.2950 1.7400 3.4150 2.7900 ;
        RECT  1.9150 1.7400 2.0350 2.7900 ;
        RECT  0.3350 1.5600 0.4550 2.7900 ;
        END
    END VDD
END NOR2X4

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3700 1.0600 1.6900 1.1800 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.3000 0.8900 1.4200 ;
        RECT  0.6500 1.3000 0.8000 1.7250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        RECT  1.0100 1.3200 1.9300 1.4400 ;
        RECT  1.8100 0.8200 1.9300 1.4400 ;
        RECT  0.5900 0.8200 1.9300 0.9400 ;
        RECT  1.4300 0.6500 1.5500 0.9400 ;
        RECT  1.0100 1.3200 1.1300 2.2100 ;
        RECT  0.5900 0.6500 0.7100 0.9400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.8500 -0.1800 1.9700 0.7000 ;
        RECT  1.0100 -0.1800 1.1300 0.7000 ;
        RECT  0.1700 -0.1800 0.2900 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.6500 1.5600 1.7700 2.7900 ;
        RECT  0.2100 1.5600 0.3300 2.7900 ;
        END
    END VDD
END NOR2X2

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.4500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 1.0000 0.8200 1.3800 ;
        RECT  0.6500 1.1750 0.8000 1.5500 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7850 0.5100 1.2350 ;
        RECT  0.3600 0.7600 0.4800 1.2350 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3196  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.9400 0.7600 1.0600 2.0050 ;
        RECT  0.6300 0.7600 1.0600 0.8800 ;
        RECT  0.6300 0.5450 0.7500 0.8800 ;
        RECT  0.6200 0.4250 0.7400 0.6650 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.4500 0.1800 ;
        RECT  1.0400 -0.1800 1.1600 0.6400 ;
        RECT  0.2000 -0.1800 0.3200 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.4500 2.7900 ;
        RECT  0.2000 1.3550 0.3200 2.7900 ;
        END
    END VDD
END NOR2X1

MACRO NOR2BXL
    CLASS CORE ;
    FOREIGN NOR2BXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0000 0.5100 1.4900 ;
        RECT  0.3600 1.0000 0.5100 1.4650 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.2350 1.3600 ;
        RECT  1.1150 1.1200 1.2350 1.3600 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1776  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 0.7600 0.6750 0.8800 ;
        RECT  0.5550 0.4000 0.6750 0.8800 ;
        RECT  0.3350 1.6100 0.4550 1.8500 ;
        RECT  0.1200 1.6100 0.4550 1.7300 ;
        RECT  0.0700 1.4650 0.2400 1.7250 ;
        RECT  0.1200 0.7600 0.2400 1.7300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.6100 1.0950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5150 1.7300 1.3950 1.7300 1.3950 1.0000 0.8150 1.0000 0.8150 0.7600 0.9350 0.7600
                 0.9350 0.8800 1.3950 0.8800 1.3950 0.4000 1.5150 0.4000 ;
    END
END NOR2BXL

MACRO NOR2BX4
    CLASS CORE ;
    FOREIGN NOR2BX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4950 1.2400 3.6150 1.4800 ;
        RECT  3.2900 1.3600 3.6150 1.4800 ;
        RECT  3.2600 1.4650 3.4100 1.7250 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2500 2.5550 1.3700 ;
        RECT  2.0450 1.2300 2.3050 1.3800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9664  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1750 0.7300 3.1950 0.8500 ;
        RECT  3.0750 0.6100 3.1950 0.8500 ;
        RECT  2.3550 1.5000 2.4750 2.2100 ;
        RECT  2.2350 0.6100 2.3550 0.8500 ;
        RECT  0.1750 1.5000 2.4750 1.6200 ;
        RECT  1.3950 0.6100 1.5150 0.8500 ;
        RECT  1.0750 1.5000 1.1950 2.2100 ;
        RECT  0.5550 0.6100 0.6750 0.8500 ;
        RECT  0.1750 1.2300 0.5650 1.3800 ;
        RECT  0.1750 0.7300 0.2950 1.6200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.4950 -0.1800 3.6150 0.8500 ;
        RECT  2.5950 0.4800 2.8350 0.6000 ;
        RECT  2.5950 -0.1800 2.7150 0.6000 ;
        RECT  1.7550 0.4800 1.9950 0.6000 ;
        RECT  1.7550 -0.1800 1.8750 0.6000 ;
        RECT  0.9150 0.4800 1.1550 0.6000 ;
        RECT  0.9150 -0.1800 1.0350 0.6000 ;
        RECT  0.0750 0.4800 0.3150 0.6000 ;
        RECT  0.0750 -0.1800 0.1950 0.6000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.2950 1.8450 3.4150 2.7900 ;
        RECT  1.7150 1.7400 1.8350 2.7900 ;
        RECT  0.3350 1.7400 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.0350 0.9900 3.8950 0.9900 3.8950 1.8000 3.7750 1.8000 3.7750 1.1100 3.3350 1.1100
                 3.3350 1.1300 3.0950 1.1300 3.0950 1.1100 1.9250 1.1100 1.9250 1.1300 1.6850 1.1300
                 1.6850 1.1100 0.4150 1.1100 0.4150 0.9900 3.7750 0.9900 3.7750 0.8700 3.9150 0.8700
                 3.9150 0.6100 4.0350 0.6100 ;
    END
END NOR2BX4

MACRO NOR2BX2
    CLASS CORE ;
    FOREIGN NOR2BX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.4650 1.3800 1.7250 ;
        RECT  1.2300 1.3400 1.3500 1.7250 ;
        RECT  1.2150 1.2200 1.3350 1.4600 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 1.2400 2.0150 1.5850 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3350 0.6900 1.5750 0.8100 ;
        RECT  0.1750 0.7400 1.4550 0.8600 ;
        RECT  0.9750 1.3200 1.0950 2.2100 ;
        RECT  0.1750 1.3200 1.0950 1.4400 ;
        RECT  0.4950 0.6900 0.7350 0.8600 ;
        RECT  0.0700 1.1750 0.2950 1.4350 ;
        RECT  0.1750 0.7400 0.2950 1.4400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8150 -0.1800 1.9350 0.8600 ;
        RECT  0.9150 0.5000 1.1550 0.6200 ;
        RECT  0.9150 -0.1800 1.0350 0.6200 ;
        RECT  0.0750 0.5000 0.3150 0.6200 ;
        RECT  0.0750 -0.1800 0.1950 0.6200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.6950 1.8450 1.8150 2.7900 ;
        RECT  0.3350 1.5600 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3550 0.9800 2.2950 0.9800 2.2950 1.8000 2.1750 1.8000 2.1750 1.1000 1.7150 1.1000
                 1.7150 1.1500 1.4750 1.1500 1.4750 1.1000 0.6550 1.1000 0.6550 1.1300 0.4150 1.1300
                 0.4150 1.0100 0.5350 1.0100 0.5350 0.9800 2.1750 0.9800 2.1750 0.8600 2.2350 0.8600
                 2.2350 0.6200 2.3550 0.6200 ;
    END
END NOR2BX2

MACRO NOR2BX1
    CLASS CORE ;
    FOREIGN NOR2BX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0000 0.5100 1.4750 ;
        RECT  0.3600 1.0000 0.5100 1.4500 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1350 1.1650 1.2550 1.4400 ;
        RECT  0.8850 1.2150 1.2550 1.3800 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3196  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.5900 0.6750 0.8500 ;
        RECT  0.1200 0.7600 0.5950 0.8800 ;
        RECT  0.4750 0.7300 0.6750 0.8500 ;
        RECT  0.2750 1.5950 0.3950 2.2100 ;
        RECT  0.1200 1.5950 0.3950 1.7150 ;
        RECT  0.1200 0.7600 0.2400 1.7150 ;
        RECT  0.0700 0.8850 0.2400 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.8050 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9150 1.5600 1.0350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5150 1.8000 1.3950 1.8000 1.3950 1.0450 1.0150 1.0450 1.0150 1.0900 0.7150 1.0900
                 0.7150 0.9700 0.8950 0.9700 0.8950 0.9250 1.3950 0.9250 1.3950 0.5650 1.5150 0.5650 ;
    END
END NOR2BX1

MACRO NAND4XL
    CLASS CORE ;
    FOREIGN NAND4XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4150 1.0250 1.5350 1.2650 ;
        RECT  1.2300 1.0250 1.5350 1.1450 ;
        RECT  1.2300 0.8850 1.3800 1.1450 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 0.8800 1.1100 1.2850 ;
        RECT  0.9400 0.7500 1.0900 1.1450 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.5950 0.8000 1.0450 ;
        RECT  0.6700 0.5950 0.7900 1.2450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.5950 0.5100 1.0150 ;
        RECT  0.3500 0.8050 0.4700 1.2450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2976  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4350 1.4050 1.7750 1.5250 ;
        RECT  1.6550 0.7850 1.7750 1.5250 ;
        RECT  1.5200 0.6650 1.6750 0.8550 ;
        RECT  1.5200 0.5950 1.6700 0.8550 ;
        RECT  1.5500 0.7850 1.7750 0.9050 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  0.1350 -0.1800 0.2550 0.3850 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.7750 1.9850 1.8950 2.7900 ;
        RECT  0.8550 1.9850 0.9750 2.7900 ;
        RECT  0.1350 1.9850 0.2550 2.7900 ;
        END
    END VDD
END NAND4XL

MACRO NAND4X8
    CLASS CORE ;
    FOREIGN NAND4X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6050 1.0300 10.9700 1.1500 ;
        RECT  9.5850 0.9400 9.8450 1.0900 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9000 1.1750 8.0500 1.4350 ;
        RECT  7.8650 1.0550 7.9850 1.2950 ;
        RECT  6.6550 1.1750 8.0500 1.2950 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7750 1.1750 5.0750 1.2950 ;
        RECT  3.8400 1.1750 3.9900 1.4350 ;
        RECT  3.7750 1.0550 3.8950 1.2950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.1750 2.0750 1.2950 ;
        RECT  1.9550 1.0550 2.0750 1.2950 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.9616  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3450 0.7000 12.1050 0.8200 ;
        RECT  11.5050 1.4700 11.6250 2.2100 ;
        RECT  0.5550 1.5550 11.6250 1.6750 ;
        RECT  11.0900 0.7000 11.2400 1.1450 ;
        RECT  11.0900 0.7000 11.2100 1.6750 ;
        RECT  10.6450 1.4700 10.7650 2.2100 ;
        RECT  9.8050 1.4650 9.9250 2.2100 ;
        RECT  8.9650 1.4700 9.0850 2.2100 ;
        RECT  8.1150 1.5550 8.2350 2.2100 ;
        RECT  7.2750 1.4650 7.3950 2.2100 ;
        RECT  6.4350 1.4650 6.5550 2.2100 ;
        RECT  5.5950 1.4700 5.7150 2.2100 ;
        RECT  4.7550 1.4700 4.8750 2.2100 ;
        RECT  3.9150 1.5550 4.0350 2.2100 ;
        RECT  3.0750 1.4700 3.1950 2.2100 ;
        RECT  2.2350 1.5550 2.3550 2.2100 ;
        RECT  1.3950 1.4650 1.5150 2.2100 ;
        RECT  0.5550 1.4650 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  2.6550 -0.1800 2.7750 0.6450 ;
        RECT  1.8150 -0.1800 1.9350 0.6450 ;
        RECT  0.9750 -0.1800 1.0950 0.6450 ;
        RECT  0.1350 -0.1800 0.2550 0.6450 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.9250 1.4700 12.0450 2.7900 ;
        RECT  11.0850 1.7950 11.2050 2.7900 ;
        RECT  10.2250 1.7950 10.3450 2.7900 ;
        RECT  9.3850 1.7950 9.5050 2.7900 ;
        RECT  8.5350 1.7950 8.6550 2.7900 ;
        RECT  7.6950 1.7950 7.8150 2.7900 ;
        RECT  6.8550 1.7950 6.9750 2.7900 ;
        RECT  6.0150 1.7950 6.1350 2.7900 ;
        RECT  5.1750 1.7950 5.2950 2.7900 ;
        RECT  4.3350 1.7950 4.4550 2.7900 ;
        RECT  3.4950 1.7950 3.6150 2.7900 ;
        RECT  2.6550 1.7950 2.7750 2.7900 ;
        RECT  1.8150 1.7950 1.9350 2.7900 ;
        RECT  0.9750 1.7950 1.0950 2.7900 ;
        RECT  0.1350 1.4650 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        RECT  6.3750 0.4600 11.6850 0.5800 ;
        POLYGON  8.7450 0.8200 6.0150 0.8200 6.0150 0.5950 3.4350 0.5950 3.4350 0.4750 6.1350 0.4750
                 6.1350 0.7000 8.7450 0.7000 ;
        POLYGON  5.7750 0.8350 5.6550 0.8350 5.6550 0.8850 0.6150 0.8850 0.6150 0.8400 0.4950 0.8400
                 0.4950 0.7200 0.7350 0.7200 0.7350 0.7650 1.3350 0.7650 1.3350 0.7150 1.5750 0.7150
                 1.5750 0.7650 2.1750 0.7650 2.1750 0.7150 2.4150 0.7150 2.4150 0.7650 3.0150 0.7650
                 3.0150 0.7150 3.2550 0.7150 3.2550 0.7650 3.8550 0.7650 3.8550 0.7150 4.0950 0.7150
                 4.0950 0.7650 4.6950 0.7650 4.6950 0.7150 4.9350 0.7150 4.9350 0.7650 5.5350 0.7650
                 5.5350 0.7150 5.7750 0.7150 ;
    END
END NAND4X8

MACRO NAND4X6
    CLASS CORE ;
    FOREIGN NAND4X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0750 1.1700 7.7350 1.2900 ;
        RECT  6.9750 1.2300 7.2350 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2900 1.1750 5.5950 1.3300 ;
        RECT  5.4750 1.0900 5.5950 1.3300 ;
        RECT  5.2900 1.1750 5.4400 1.4350 ;
        RECT  5.0950 1.1500 5.3350 1.2700 ;
        RECT  5.2150 1.1750 5.5950 1.2950 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2950 1.1700 3.5350 1.2900 ;
        RECT  2.9700 1.1750 3.4150 1.2950 ;
        RECT  2.9700 1.1750 3.1200 1.4350 ;
        RECT  2.9950 1.1100 3.1150 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        RECT  1.2550 1.1100 1.3750 1.4350 ;
        RECT  0.9550 1.1750 1.3800 1.2950 ;
        RECT  0.8350 1.1700 1.0750 1.2900 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.9712  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9950 0.9300 8.8550 1.0500 ;
        RECT  8.7350 0.4000 8.8550 1.0500 ;
        RECT  8.2550 1.4300 8.3750 2.2100 ;
        RECT  0.6950 1.5550 8.3750 1.6750 ;
        RECT  7.9000 1.1750 8.0500 1.4350 ;
        RECT  7.9000 0.9300 8.0200 1.6750 ;
        RECT  7.8350 0.6000 7.9550 1.0500 ;
        RECT  7.4150 1.4300 7.5350 2.2100 ;
        RECT  6.9950 0.6000 7.1150 1.0500 ;
        RECT  6.5750 1.4300 6.6950 2.2100 ;
        RECT  5.7350 1.4300 5.8550 2.2100 ;
        RECT  4.8950 1.4300 5.0150 2.2100 ;
        RECT  4.0550 1.4300 4.1750 2.2100 ;
        RECT  3.2150 1.5550 3.3350 2.2100 ;
        RECT  2.3750 1.4300 2.4950 2.2100 ;
        RECT  1.5350 1.4300 1.6550 2.2100 ;
        RECT  0.6950 1.4300 0.8150 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  1.8750 -0.1800 1.9950 0.7500 ;
        RECT  1.0350 -0.1800 1.1550 0.7500 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.6750 1.4300 8.7950 2.7900 ;
        RECT  7.8350 1.7950 7.9550 2.7900 ;
        RECT  6.9950 1.7950 7.1150 2.7900 ;
        RECT  6.1550 1.7950 6.2750 2.7900 ;
        RECT  5.3150 1.7950 5.4350 2.7900 ;
        RECT  4.4750 1.7950 4.5950 2.7900 ;
        RECT  3.6350 1.7950 3.7550 2.7900 ;
        RECT  2.7950 1.7950 2.9150 2.7900 ;
        RECT  1.9550 1.7950 2.0750 2.7900 ;
        RECT  1.1150 1.7950 1.2350 2.7900 ;
        RECT  0.2750 1.4300 0.3950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.4350 0.8100 8.3150 0.8100 8.3150 0.4800 7.5350 0.4800 7.5350 0.8100 7.4150 0.8100
                 7.4150 0.4800 6.6950 0.4800 6.6950 0.9200 6.5750 0.9200 6.5750 0.4800 5.8550 0.4800
                 5.8550 0.7300 5.7350 0.7300 5.7350 0.4800 4.9550 0.4800 4.9550 0.7300 4.8350 0.7300
                 4.8350 0.3600 8.4350 0.3600 ;
        POLYGON  6.2750 0.9700 4.4150 0.9700 4.4150 0.4800 3.6750 0.4800 3.6750 0.7500 3.5550 0.7500
                 3.5550 0.4800 2.8350 0.4800 2.8350 0.7500 2.7150 0.7500 2.7150 0.3600 4.5350 0.3600
                 4.5350 0.8500 5.3150 0.8500 5.3150 0.6000 5.4350 0.6000 5.4350 0.8500 6.1550 0.8500
                 6.1550 0.6000 6.2750 0.6000 ;
        POLYGON  4.1150 0.9900 0.5550 0.9900 0.5550 0.4000 0.6750 0.4000 0.6750 0.8700 1.4550 0.8700
                 1.4550 0.4000 1.5750 0.4000 1.5750 0.8700 2.2950 0.8700 2.2950 0.4000 2.4150 0.4000
                 2.4150 0.8700 3.1350 0.8700 3.1350 0.6000 3.2550 0.6000 3.2550 0.8700 3.9950 0.8700
                 3.9950 0.6000 4.1150 0.6000 ;
    END
END NAND4X6

MACRO NAND4X4
    CLASS CORE ;
    FOREIGN NAND4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5850 1.0800 6.8250 1.2000 ;
        RECT  5.8650 1.2600 6.7050 1.3800 ;
        RECT  6.5850 1.0800 6.7050 1.3800 ;
        RECT  6.1050 1.2300 6.3650 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5050 1.0800 5.7450 1.2000 ;
        RECT  4.1350 1.2600 5.6250 1.3800 ;
        RECT  5.5050 1.0800 5.6250 1.3800 ;
        RECT  5.2350 1.2300 5.6250 1.3800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4550 1.2600 3.0350 1.3800 ;
        RECT  2.6250 1.2300 2.8850 1.3800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 1.2600 1.3150 1.3800 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.9392  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2650 0.8400 7.0250 0.9600 ;
        RECT  6.9050 0.6400 7.0250 0.9600 ;
        RECT  6.4350 1.5000 6.5550 2.2100 ;
        RECT  0.5550 1.5000 6.5550 1.6200 ;
        RECT  6.0650 0.6400 6.1850 0.9600 ;
        RECT  5.5950 1.5000 5.7150 2.2100 ;
        RECT  2.2150 0.9900 5.3850 1.1100 ;
        RECT  5.2650 0.8400 5.3850 1.1100 ;
        RECT  4.7550 1.5000 4.8750 2.2100 ;
        RECT  3.9150 1.5000 4.0350 2.2100 ;
        RECT  3.0750 1.5000 3.1950 2.2100 ;
        RECT  2.2350 1.5000 2.3550 2.2100 ;
        RECT  2.1000 1.4650 2.3350 1.7250 ;
        RECT  2.2150 0.9900 2.3350 1.7250 ;
        RECT  1.3950 1.5000 1.5150 2.2100 ;
        RECT  0.5550 1.5000 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  1.3950 -0.1800 1.5150 0.6900 ;
        RECT  0.5550 -0.1800 0.6750 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  6.8550 1.5600 6.9750 2.7900 ;
        RECT  6.0150 1.7400 6.1350 2.7900 ;
        RECT  5.1750 1.7400 5.2950 2.7900 ;
        RECT  4.3350 1.7400 4.4550 2.7900 ;
        RECT  3.4950 1.7400 3.6150 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.4450 0.6900 7.3250 0.6900 7.3250 0.4800 6.6050 0.4800 6.6050 0.6900 6.4850 0.6900
                 6.4850 0.4800 5.7650 0.4800 5.7650 0.6900 5.6450 0.6900 5.6450 0.4800 4.9050 0.4800
                 4.9050 0.6300 4.6650 0.6300 4.6650 0.4800 4.0650 0.4800 4.0650 0.6300 3.8250 0.6300
                 3.8250 0.5100 3.9450 0.5100 3.9450 0.3600 7.4450 0.3600 ;
        POLYGON  5.4050 0.7200 5.1450 0.7200 5.1450 0.8700 2.3550 0.8700 2.3550 0.8200 2.1750 0.8200
                 2.1750 0.7000 2.4750 0.7000 2.4750 0.7500 3.0750 0.7500 3.0750 0.6300 3.1950 0.6300
                 3.1950 0.7500 4.3050 0.7500 4.3050 0.6300 4.4250 0.6300 4.4250 0.7500 5.0250 0.7500
                 5.0250 0.6000 5.4050 0.6000 ;
        POLYGON  3.6750 0.6300 3.4350 0.6300 3.4350 0.5100 2.8350 0.5100 2.8350 0.6300 2.5950 0.6300
                 2.5950 0.5100 1.9350 0.5100 1.9350 0.9300 0.1350 0.9300 0.1350 0.6400 0.2550 0.6400
                 0.2550 0.8100 0.9750 0.8100 0.9750 0.6400 1.0950 0.6400 1.0950 0.8100 1.8150 0.8100
                 1.8150 0.3900 3.5550 0.3900 3.5550 0.5100 3.6750 0.5100 ;
    END
END NAND4X4

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8400 0.9700 2.0800 1.0900 ;
        RECT  1.8400 0.5950 1.9600 1.0900 ;
        RECT  1.8100 0.5950 1.9600 0.8550 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9400 2.8850 1.0900 ;
        RECT  1.3800 1.2100 2.8400 1.3300 ;
        RECT  2.7200 0.9400 2.8400 1.3300 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9600 1.4500 3.3800 1.5700 ;
        RECT  3.2600 1.2200 3.3800 1.5700 ;
        RECT  0.9600 1.1750 1.0900 1.5700 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.8400 1.2800 1.0900 1.4000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5800 1.6900 3.7000 1.8100 ;
        RECT  3.5800 1.2200 3.7000 1.8100 ;
        RECT  3.5500 1.4650 3.7000 1.8100 ;
        RECT  0.5800 1.2200 0.7000 1.8100 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9696  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8200 1.7550 3.9900 2.0150 ;
        RECT  0.6400 1.9300 3.9400 2.0500 ;
        RECT  3.8200 0.7000 3.9400 2.0500 ;
        RECT  2.2400 0.7000 3.9400 0.8200 ;
        RECT  3.5200 1.9300 3.6400 2.2100 ;
        RECT  2.5600 1.9300 2.6800 2.2100 ;
        RECT  2.1200 0.6500 2.3600 0.7700 ;
        RECT  1.6000 1.9300 1.7200 2.2100 ;
        RECT  0.6400 1.9300 0.7600 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.6800 0.4600 3.9200 0.5800 ;
        RECT  3.6800 -0.1800 3.8000 0.5800 ;
        RECT  0.4200 -0.1800 0.5400 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.9400 2.1700 4.1800 2.2900 ;
        RECT  3.9400 2.1700 4.0600 2.7900 ;
        RECT  2.9800 2.1700 3.2200 2.2900 ;
        RECT  2.9800 2.1700 3.1000 2.7900 ;
        RECT  2.0200 2.1700 2.2600 2.2900 ;
        RECT  2.0200 2.1700 2.1400 2.7900 ;
        RECT  1.0600 2.1700 1.3000 2.2900 ;
        RECT  1.0600 2.1700 1.1800 2.7900 ;
        RECT  0.2200 1.5600 0.3400 2.7900 ;
        END
    END VDD
END NAND4X2

MACRO NAND4X1
    CLASS CORE ;
    FOREIGN NAND4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 0.5950 1.6700 1.1800 ;
        RECT  1.5200 0.5950 1.6700 1.0200 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.5950 1.3800 1.0000 ;
        RECT  1.2100 0.7800 1.3300 1.2000 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8900 0.9600 1.0100 1.2000 ;
        RECT  0.6500 0.9600 1.0100 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2750 0.8850 0.5300 1.1450 ;
        RECT  0.2350 0.9400 0.4700 1.1800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5364  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7900 1.1750 1.9600 1.4350 ;
        RECT  0.6300 1.3200 1.9100 1.4400 ;
        RECT  1.7900 0.6200 1.9100 1.4400 ;
        RECT  1.4700 1.3200 1.5900 2.2100 ;
        RECT  0.6300 1.3200 0.7500 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  0.4100 -0.1800 0.5300 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.8900 1.5600 2.0100 2.7900 ;
        RECT  1.0500 1.5600 1.1700 2.7900 ;
        RECT  0.2100 1.5600 0.3300 2.7900 ;
        END
    END VDD
END NAND4X1

MACRO NAND4BXL
    CLASS CORE ;
    FOREIGN NAND4BXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.8500 0.5100 1.3500 ;
        RECT  0.3600 0.8500 0.5100 1.3200 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.9050 0.9350 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.8850 1.3800 1.2750 ;
        RECT  1.1400 0.8300 1.2600 1.2300 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7200 1.1750 2.0150 1.4450 ;
        RECT  1.7200 1.1750 1.9600 1.4600 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2976  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3350 1.6500 1.5750 1.7700 ;
        RECT  1.3350 1.4700 1.4550 1.7700 ;
        RECT  0.1200 1.4700 1.4550 1.5900 ;
        RECT  0.4950 1.4700 0.7350 1.7700 ;
        RECT  0.0700 0.5950 0.4550 0.7300 ;
        RECT  0.3350 0.4900 0.4550 0.7300 ;
        RECT  0.1200 0.5950 0.2400 1.5900 ;
        RECT  0.0700 0.5950 0.2400 0.8550 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.6200 -0.1800 1.7400 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8750 2.2300 1.9950 2.7900 ;
        RECT  0.9150 2.2300 1.0350 2.7900 ;
        RECT  0.1350 1.7100 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4750 1.8300 2.3550 1.8300 2.3550 1.7100 2.1350 1.7100 2.1350 1.0100 1.5000 1.0100
                 1.5000 0.8900 2.1350 0.8900 2.1350 0.7300 2.0400 0.7300 2.0400 0.4900 2.1600 0.4900
                 2.1600 0.6100 2.2550 0.6100 2.2550 1.5900 2.4750 1.5900 ;
    END
END NAND4BXL

MACRO NAND4BX4
    CLASS CORE ;
    FOREIGN NAND4BX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0350 1.0800 7.6350 1.2000 ;
        RECT  7.0350 1.0800 7.2750 1.3500 ;
        RECT  6.6750 1.2600 7.2350 1.3800 ;
        RECT  6.9750 1.2300 7.2750 1.3500 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3150 1.0800 6.5550 1.2000 ;
        RECT  4.9450 1.2600 6.4350 1.3800 ;
        RECT  6.3150 1.0800 6.4350 1.3800 ;
        RECT  6.1050 1.2300 6.4350 1.3800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2650 1.2600 3.8450 1.3800 ;
        RECT  3.4950 1.2300 3.7550 1.3800 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2750 1.0000 0.3950 1.2400 ;
        RECT  0.0700 1.0000 0.3950 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.9392  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0750 0.8400 7.8350 0.9600 ;
        RECT  7.7150 0.6400 7.8350 0.9600 ;
        RECT  7.2450 1.5000 7.3650 2.2100 ;
        RECT  1.3650 1.5000 7.3650 1.6200 ;
        RECT  6.8750 0.6400 6.9950 0.9600 ;
        RECT  6.4050 1.5000 6.5250 2.2100 ;
        RECT  3.0250 0.9900 6.1950 1.1100 ;
        RECT  6.0750 0.8400 6.1950 1.1100 ;
        RECT  5.5650 1.5000 5.6850 2.2100 ;
        RECT  4.7250 1.5000 4.8450 2.2100 ;
        RECT  3.8850 1.5000 4.0050 2.2100 ;
        RECT  3.0450 1.5000 3.1650 2.2100 ;
        RECT  2.9700 1.4650 3.1450 1.7250 ;
        RECT  3.0250 0.9900 3.1450 1.7250 ;
        RECT  2.2050 1.5000 2.3250 2.2100 ;
        RECT  1.3650 1.5000 1.4850 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  2.2050 -0.1800 2.3250 0.6900 ;
        RECT  1.3650 -0.1800 1.4850 0.6900 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.6650 1.5600 7.7850 2.7900 ;
        RECT  6.8250 1.7400 6.9450 2.7900 ;
        RECT  5.9850 1.7400 6.1050 2.7900 ;
        RECT  5.1450 1.7400 5.2650 2.7900 ;
        RECT  4.3050 1.7400 4.4250 2.7900 ;
        RECT  3.4650 1.7400 3.5850 2.7900 ;
        RECT  2.6250 1.7400 2.7450 2.7900 ;
        RECT  1.7850 1.7400 1.9050 2.7900 ;
        RECT  0.9450 1.5600 1.0650 2.7900 ;
        RECT  0.1350 1.3600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2550 0.6900 8.1350 0.6900 8.1350 0.4800 7.4150 0.4800 7.4150 0.6900 7.2950 0.6900
                 7.2950 0.4800 6.5750 0.4800 6.5750 0.6900 6.4550 0.6900 6.4550 0.4800 5.7150 0.4800
                 5.7150 0.6300 5.4750 0.6300 5.4750 0.4800 4.8750 0.4800 4.8750 0.6300 4.6350 0.6300
                 4.6350 0.5100 4.7550 0.5100 4.7550 0.3600 8.2550 0.3600 ;
        POLYGON  6.2150 0.7200 5.9550 0.7200 5.9550 0.8700 3.1650 0.8700 3.1650 0.8200 2.9850 0.8200
                 2.9850 0.7000 3.2850 0.7000 3.2850 0.7500 3.8850 0.7500 3.8850 0.6300 4.0050 0.6300
                 4.0050 0.7500 5.1150 0.7500 5.1150 0.6300 5.2350 0.6300 5.2350 0.7500 5.8350 0.7500
                 5.8350 0.6000 6.2150 0.6000 ;
        POLYGON  4.4850 0.6300 4.2450 0.6300 4.2450 0.5100 3.6450 0.5100 3.6450 0.6300 3.4050 0.6300
                 3.4050 0.5100 2.7450 0.5100 2.7450 0.9300 0.9450 0.9300 0.9450 0.6400 1.0650 0.6400
                 1.0650 0.8100 1.7850 0.8100 1.7850 0.6400 1.9050 0.6400 1.9050 0.8100 2.6250 0.8100
                 2.6250 0.3900 4.3650 0.3900 4.3650 0.5100 4.4850 0.5100 ;
        POLYGON  2.1250 1.3600 0.6750 1.3600 0.6750 2.0100 0.5550 2.0100 0.5550 0.6800 0.6750 0.6800
                 0.6750 1.2400 2.1250 1.2400 ;
    END
END NAND4BX4

MACRO NAND4BX2
    CLASS CORE ;
    FOREIGN NAND4BX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0350 1.2100 4.3350 1.4400 ;
        RECT  4.0750 1.1850 4.3350 1.4400 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 1.2600 3.3150 1.4350 ;
        RECT  2.9150 1.2300 3.1750 1.4350 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.1800 2.5950 1.4500 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2950 1.2200 0.5650 1.3800 ;
        RECT  0.1750 1.1200 0.4150 1.2500 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9696  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1950 0.6500 4.4350 0.7700 ;
        RECT  2.0950 0.9400 4.3150 1.0600 ;
        RECT  4.1950 0.6500 4.3150 1.0600 ;
        RECT  3.9350 1.5600 4.0550 2.2100 ;
        RECT  1.4150 1.5700 4.0550 1.6900 ;
        RECT  3.0950 1.5600 3.2150 2.2100 ;
        RECT  2.2550 1.5700 2.3750 2.2100 ;
        RECT  2.1000 1.5700 2.3750 2.0150 ;
        RECT  2.0950 0.9400 2.2150 1.6900 ;
        RECT  1.4150 1.5600 1.5350 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  1.3450 -0.1800 1.4650 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  4.3550 1.5600 4.4750 2.7900 ;
        RECT  3.5150 1.8100 3.6350 2.7900 ;
        RECT  2.6750 1.8100 2.7950 2.7900 ;
        RECT  1.8350 1.8100 1.9550 2.7900 ;
        RECT  0.9950 1.7700 1.1150 2.7900 ;
        RECT  0.2650 1.5000 0.3850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.7950 0.6500 4.6750 0.6500 4.6750 0.5300 3.9550 0.5300 3.9550 0.6500 3.8350 0.6500
                 3.8350 0.5300 3.1750 0.5300 3.1750 0.5800 2.9350 0.5800 2.9350 0.4600 3.0550 0.4600
                 3.0550 0.4100 4.7950 0.4100 ;
        POLYGON  3.5950 0.7700 3.4750 0.7700 3.4750 0.8200 2.2450 0.8200 2.2450 0.7700 2.1250 0.7700
                 2.1250 0.6500 2.3650 0.6500 2.3650 0.7000 3.3550 0.7000 3.3550 0.6500 3.5950 0.6500 ;
        POLYGON  2.7850 0.5800 2.5450 0.5800 2.5450 0.5300 1.8850 0.5300 1.8850 0.8800 0.9250 0.8800
                 0.9250 0.5900 1.0450 0.5900 1.0450 0.7600 1.7650 0.7600 1.7650 0.4100 2.6650 0.4100
                 2.6650 0.4600 2.7850 0.4600 ;
        POLYGON  1.3350 1.3200 0.8050 1.3200 0.8050 1.6200 0.6850 1.6200 0.6850 1.1000 0.5350 1.1000
                 0.5350 0.6800 0.6550 0.6800 0.6550 0.9800 0.8050 0.9800 0.8050 1.2000 1.3350 1.2000 ;
    END
END NAND4BX2

MACRO NAND4BX1
    CLASS CORE ;
    FOREIGN NAND4BX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7850 0.5100 1.2400 ;
        RECT  0.3900 0.7600 0.5100 1.2400 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8900 0.9300 1.0100 1.1700 ;
        RECT  0.6500 0.9300 1.0100 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.8850 1.4150 1.2150 ;
        RECT  1.2100 0.8450 1.3650 1.1700 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0000 2.2500 1.4700 ;
        RECT  2.1000 1.0000 2.2200 1.5000 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5364  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4700 1.3600 1.5900 2.2100 ;
        RECT  0.1200 1.3600 1.5900 1.4800 ;
        RECT  0.6300 1.3600 0.7500 2.2100 ;
        RECT  0.1200 0.5200 0.5300 0.6400 ;
        RECT  0.4100 0.4000 0.5300 0.6400 ;
        RECT  0.0700 1.1750 0.2400 1.4350 ;
        RECT  0.1200 0.5200 0.2400 1.4800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.6900 -0.1800 1.8100 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.8900 1.6200 2.0100 2.7900 ;
        RECT  1.0500 1.6000 1.1700 2.7900 ;
        RECT  0.2100 1.6000 0.3300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4900 1.8000 2.3700 1.8000 2.3700 0.8800 1.9800 0.8800 1.9800 1.1100 1.6300 1.1100
                 1.6300 0.9900 1.8600 0.9900 1.8600 0.7600 2.1700 0.7600 2.1700 0.5900 2.2900 0.5900
                 2.2900 0.7100 2.4900 0.7100 ;
    END
END NAND4BX1

MACRO NAND4BBXL
    CLASS CORE ;
    FOREIGN NAND4BBXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2750 0.9400 0.3950 1.1800 ;
        RECT  0.0700 0.9400 0.3950 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4250 1.3200 2.6650 1.5050 ;
        RECT  2.3350 1.2300 2.5950 1.4400 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.1750 1.6700 1.5200 ;
        RECT  1.4250 1.3250 1.5450 1.6700 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2300 1.1450 1.5000 ;
        RECT  0.8150 1.3600 1.0550 1.6100 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2976  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9450 0.6950 2.0650 2.0900 ;
        RECT  1.1050 1.7900 2.0650 1.9100 ;
        RECT  1.8100 1.4650 2.0650 1.9100 ;
        RECT  1.0050 0.6950 2.0650 0.8150 ;
        RECT  1.1050 1.7900 1.2250 2.0900 ;
        RECT  0.8850 0.5950 1.1250 0.7150 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.3250 -0.1800 2.4450 0.7750 ;
        RECT  0.1350 -0.1800 0.2550 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3650 1.9700 2.4850 2.7900 ;
        RECT  1.4650 2.0300 1.7050 2.1500 ;
        RECT  1.4650 2.0300 1.5850 2.7900 ;
        RECT  0.6850 1.9700 0.8050 2.7900 ;
        RECT  0.1350 1.4600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.9250 0.7150 2.9050 0.7150 2.9050 2.0900 2.7850 2.0900 2.7850 1.1100 2.1850 1.1100
                 2.1850 0.9900 2.7850 0.9900 2.7850 0.7150 2.6850 0.7150 2.6850 0.5950 2.9250 0.5950 ;
        POLYGON  1.8250 1.0550 0.6750 1.0550 0.6750 1.5800 0.5550 1.5800 0.5550 0.5250 0.6750 0.5250
                 0.6750 0.9350 1.8250 0.9350 ;
    END
END NAND4BBXL

MACRO NAND4BBX4
    CLASS CORE ;
    FOREIGN NAND4BBX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0100 0.5100 1.4650 ;
        RECT  0.3750 1.0100 0.4950 1.4950 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0200 0.8350 1.3900 ;
        RECT  0.6500 1.0700 0.8000 1.4350 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5450 1.0300 5.7300 1.4350 ;
        RECT  5.5450 1.0150 5.6650 1.4350 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0850 0.9500 7.2050 1.4000 ;
        RECT  7.0300 0.7750 7.1800 1.2050 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.9392  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2050 0.6050 8.3250 0.8450 ;
        RECT  8.0250 0.7250 8.3250 0.8450 ;
        RECT  7.3650 0.7750 8.1450 0.8950 ;
        RECT  7.9550 1.5600 8.0750 2.2100 ;
        RECT  7.7750 1.5600 8.0750 1.6800 ;
        RECT  2.0450 1.5550 7.8950 1.6700 ;
        RECT  7.7750 0.7750 7.8950 1.6800 ;
        RECT  2.0750 1.5600 8.0750 1.6750 ;
        RECT  7.3650 0.6050 7.4850 0.8950 ;
        RECT  7.1150 1.5550 7.2350 2.2100 ;
        RECT  6.2750 1.5550 6.3950 2.2100 ;
        RECT  5.4350 1.5550 5.5550 2.2100 ;
        RECT  4.5950 1.5550 4.7150 2.2100 ;
        RECT  3.7550 1.5550 3.8750 2.2100 ;
        RECT  2.9150 1.5550 3.0350 2.2100 ;
        RECT  2.0450 1.5200 2.3050 1.6700 ;
        RECT  2.0750 1.5200 2.1950 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  2.7150 0.4750 2.9550 0.5950 ;
        RECT  2.8350 -0.1800 2.9550 0.5950 ;
        RECT  1.8750 0.4750 2.1150 0.5950 ;
        RECT  1.8750 -0.1800 1.9950 0.5950 ;
        RECT  0.5550 -0.1800 0.6750 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.3750 1.5600 8.4950 2.7900 ;
        RECT  7.5350 1.7950 7.6550 2.7900 ;
        RECT  6.6950 1.7950 6.8150 2.7900 ;
        RECT  5.8550 1.7950 5.9750 2.7900 ;
        RECT  5.0150 1.7950 5.1350 2.7900 ;
        RECT  4.1750 1.7950 4.2950 2.7900 ;
        RECT  3.3350 1.7950 3.4550 2.7900 ;
        RECT  2.4950 1.7950 2.6150 2.7900 ;
        RECT  1.6550 1.5600 1.7750 2.7900 ;
        RECT  0.5550 1.6150 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.7450 0.6550 8.6250 0.6550 8.6250 0.4850 7.9050 0.4850 7.9050 0.6550 7.7850 0.6550
                 7.7850 0.4850 7.0650 0.4850 7.0650 0.6550 6.9450 0.6550 6.9450 0.4850 6.2250 0.4850
                 6.2250 0.6550 6.1050 0.6550 6.1050 0.4850 5.3850 0.4850 5.3850 0.6550 5.2650 0.6550
                 5.2650 0.3650 8.7450 0.3650 ;
        POLYGON  6.6450 0.8950 3.7950 0.8950 3.7950 0.8850 3.6150 0.8850 3.6150 0.6050 3.7350 0.6050
                 3.7350 0.7650 3.9150 0.7650 3.9150 0.7750 4.4550 0.7750 4.4550 0.6050 4.5750 0.6050
                 4.5750 0.7750 5.6850 0.7750 5.6850 0.6050 5.8050 0.6050 5.8050 0.7750 6.5250 0.7750
                 6.5250 0.6050 6.6450 0.6050 ;
        POLYGON  4.9950 0.6550 4.8750 0.6550 4.8750 0.4850 4.1550 0.4850 4.1550 0.6550 4.0350 0.6550
                 4.0350 0.4850 3.3750 0.4850 3.3750 0.5950 3.2700 0.5950 3.2700 0.8350 2.4750 0.8350
                 2.4750 0.8450 2.3550 0.8450 2.3550 0.8350 1.6350 0.8350 1.6350 0.8450 1.5150 0.8450
                 1.5150 0.6050 1.6350 0.6050 1.6350 0.7150 2.3550 0.7150 2.3550 0.6050 2.4750 0.6050
                 2.4750 0.7150 3.1500 0.7150 3.1500 0.5950 3.1350 0.5950 3.1350 0.4750 3.2400 0.4750
                 3.2400 0.3650 4.9950 0.3650 ;
        POLYGON  3.6750 1.1250 1.2750 1.1250 1.2750 0.4800 0.9150 0.4800 0.9150 0.8900 0.2400 0.8900
                 0.2400 1.5850 0.2550 1.5850 0.2550 2.2100 0.1350 2.2100 0.1350 1.7050 0.1200 1.7050
                 0.1200 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000 0.2550 0.7700 0.7950 0.7700
                 0.7950 0.3600 1.3950 0.3600 1.3950 1.0050 3.6750 1.0050 ;
        POLYGON  1.9750 1.4000 1.1550 1.4000 1.1550 1.5200 1.0950 1.5200 1.0950 2.2100 0.9750 2.2100
                 0.9750 1.4000 1.0350 1.4000 1.0350 0.6000 1.1550 0.6000 1.1550 1.2800 1.9750 1.2800 ;
    END
END NAND4BBX4

MACRO NAND4BBX2
    CLASS CORE ;
    FOREIGN NAND4BBX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.8000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4450 1.1800 0.5650 1.6700 ;
        RECT  0.3050 1.1800 0.5650 1.4000 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.5200 1.1450 1.7050 ;
        RECT  0.8850 1.3300 1.0050 1.7050 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0950 1.0300 4.2800 1.4350 ;
        RECT  4.0950 1.0150 4.2150 1.4350 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8150 1.0750 4.9350 1.3800 ;
        RECT  4.7100 0.8800 4.8600 1.1950 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9696  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0750 0.6050 5.1950 0.8450 ;
        RECT  4.8750 1.5550 5.1750 1.6800 ;
        RECT  5.0550 0.7250 5.1750 1.6800 ;
        RECT  4.8750 1.5550 4.9950 2.2100 ;
        RECT  2.3550 1.5550 5.1750 1.6750 ;
        RECT  4.0350 1.5550 4.1550 2.2100 ;
        RECT  3.1950 1.5550 3.3150 2.2100 ;
        RECT  2.3350 1.5200 2.5950 1.6700 ;
        RECT  2.3550 1.5200 2.4750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.8000 0.1800 ;
        RECT  2.1050 0.4750 2.3450 0.5950 ;
        RECT  2.2250 -0.1800 2.3450 0.5950 ;
        RECT  0.6850 -0.1800 0.8050 0.8200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.8000 2.7900 ;
        RECT  5.2950 1.5600 5.4150 2.7900 ;
        RECT  4.4550 1.7950 4.5750 2.7900 ;
        RECT  3.6150 1.7950 3.7350 2.7900 ;
        RECT  2.7750 1.7950 2.8950 2.7900 ;
        RECT  1.9350 1.5600 2.0550 2.7900 ;
        RECT  0.6250 1.8250 0.7450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.6150 0.6550 5.4950 0.6550 5.4950 0.4850 4.7750 0.4850 4.7750 0.6550 4.6550 0.6550
                 4.6550 0.4850 3.9350 0.4850 3.9350 0.6550 3.8150 0.6550 3.8150 0.3650 5.6150 0.3650 ;
        POLYGON  4.3550 0.8950 3.1850 0.8950 3.1850 0.8850 3.0050 0.8850 3.0050 0.6050 3.1250 0.6050
                 3.1250 0.7650 3.3050 0.7650 3.3050 0.7750 4.2350 0.7750 4.2350 0.6050 4.3550 0.6050 ;
        POLYGON  3.5450 0.6550 3.4250 0.6550 3.4250 0.4850 2.7650 0.4850 2.7650 0.5950 2.6600 0.5950
                 2.6600 0.8350 1.8650 0.8350 1.8650 0.8450 1.7450 0.8450 1.7450 0.6050 1.8650 0.6050
                 1.8650 0.7150 2.5400 0.7150 2.5400 0.5950 2.5250 0.5950 2.5250 0.4750 2.6300 0.4750
                 2.6300 0.3650 3.5450 0.3650 ;
        POLYGON  3.0650 1.1250 1.5050 1.1250 1.5050 0.4800 1.0450 0.4800 1.0450 1.0600 0.1850 1.0600
                 0.1850 1.7050 0.3250 1.7050 0.3250 1.9450 0.2050 1.9450 0.2050 1.8250 0.0650 1.8250
                 0.0650 0.7200 0.2050 0.7200 0.2050 0.6000 0.3250 0.6000 0.3250 0.9400 0.9250 0.9400
                 0.9250 0.3600 1.6250 0.3600 1.6250 1.0050 3.0650 1.0050 ;
        POLYGON  2.2750 1.3650 1.3850 1.3650 1.3850 1.9450 1.1650 1.9450 1.1650 2.0650 1.0450 2.0650
                 1.0450 1.8250 1.2650 1.8250 1.2650 0.8400 1.1650 0.8400 1.1650 0.6000 1.2850 0.6000
                 1.2850 0.7200 1.3850 0.7200 1.3850 1.2450 2.2750 1.2450 ;
    END
END NAND4BBX2

MACRO NAND4BBX1
    CLASS CORE ;
    FOREIGN NAND4BBX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1600 0.9250 0.4000 1.1650 ;
        RECT  0.0600 0.8850 0.3200 1.1450 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7700 1.1300 2.9100 1.4400 ;
        RECT  2.6250 1.2300 2.9100 1.4150 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5100 0.9900 1.6700 1.4350 ;
        RECT  1.5100 0.9650 1.6350 1.4350 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9700 1.2000 1.2100 1.3900 ;
        RECT  0.8850 1.2300 1.1450 1.4450 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5364  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2900 1.5550 2.2700 1.6750 ;
        RECT  2.1500 0.4850 2.2700 1.6750 ;
        RECT  2.1300 1.4650 2.2500 2.2100 ;
        RECT  0.9700 0.4850 2.2700 0.6050 ;
        RECT  2.1000 1.4650 2.2500 1.7250 ;
        RECT  1.2900 1.5550 1.4100 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.3900 -0.1800 2.5100 0.6600 ;
        RECT  0.1400 -0.1800 0.2600 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.5500 1.5600 2.6700 2.7900 ;
        RECT  1.7100 1.7950 1.8300 2.7900 ;
        RECT  0.8700 1.7300 0.9900 2.7900 ;
        RECT  0.1400 1.4600 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1500 1.8000 3.0300 1.8000 3.0300 1.0100 2.6500 1.0100 2.6500 1.1100 2.3900 1.1100
                 2.3900 0.9900 2.5300 0.9900 2.5300 0.8900 2.9500 0.8900 2.9500 0.6100 3.0700 0.6100
                 3.0700 0.7700 3.1500 0.7700 ;
        POLYGON  2.0300 1.1100 1.7900 1.1100 1.7900 0.8450 0.6800 0.8450 0.6800 1.5800 0.5600 1.5800
                 0.5600 0.5250 0.6800 0.5250 0.6800 0.7250 1.9100 0.7250 1.9100 0.9900 2.0300 0.9900 ;
    END
END NAND4BBX1

MACRO NAND3XL
    CLASS CORE ;
    FOREIGN NAND3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6950 1.0550 0.8150 1.4850 ;
        RECT  0.6500 0.8850 0.8000 1.3000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3550 1.0600 0.5100 1.5150 ;
        RECT  0.3550 1.0400 0.4750 1.5150 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0250 1.0250 1.1750 1.2650 ;
        RECT  0.9400 0.8850 1.1150 1.1450 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4850 1.6050 1.6050 1.8450 ;
        RECT  0.6300 1.6050 1.6050 1.7250 ;
        RECT  1.2300 1.4650 1.4150 1.7250 ;
        RECT  1.2950 0.6800 1.4150 1.7250 ;
        RECT  0.4950 1.6350 0.7500 1.7550 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.1950 -0.1800 0.3150 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.0050 2.1550 1.1250 2.7900 ;
        RECT  0.1350 1.6350 0.2550 2.7900 ;
        END
    END VDD
END NAND3XL

MACRO NAND3X8
    CLASS CORE ;
    FOREIGN NAND3X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5550 1.0500 8.7950 1.1700 ;
        RECT  8.5550 0.7300 8.6750 1.1700 ;
        RECT  5.6400 0.7300 8.6750 0.8500 ;
        RECT  6.3150 1.0300 6.5550 1.1500 ;
        RECT  6.4350 0.7300 6.5550 1.1500 ;
        RECT  1.5500 0.7250 5.7600 0.8450 ;
        RECT  4.0500 1.0300 4.2900 1.1500 ;
        RECT  4.0500 0.7250 4.1700 1.1500 ;
        RECT  1.4300 1.0350 1.6700 1.1550 ;
        RECT  1.5500 0.7250 1.6700 1.1550 ;
        RECT  1.5200 0.8850 1.6700 1.1550 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7650 1.0300 8.4350 1.1500 ;
        RECT  8.1350 1.0300 8.3950 1.3800 ;
        RECT  6.9700 0.9700 7.8850 1.0900 ;
        RECT  6.7050 1.0500 7.1950 1.1700 ;
        RECT  5.9100 1.2700 6.8250 1.3900 ;
        RECT  6.7050 1.0500 6.8250 1.3900 ;
        RECT  5.9100 1.1100 6.0300 1.3900 ;
        RECT  5.3800 1.1100 6.0300 1.2300 ;
        RECT  5.3800 0.9650 5.5000 1.2300 ;
        RECT  4.7800 0.9650 5.5000 1.0850 ;
        RECT  4.4100 1.1050 4.9000 1.2250 ;
        RECT  4.7800 0.9650 4.9000 1.2250 ;
        RECT  3.8100 1.2700 4.5300 1.3900 ;
        RECT  4.4100 1.1050 4.5300 1.3900 ;
        RECT  3.8100 1.0500 3.9300 1.3900 ;
        RECT  3.0150 1.0500 3.9300 1.1700 ;
        RECT  2.2200 0.9650 3.1350 1.0850 ;
        RECT  1.9350 1.0450 2.3400 1.1650 ;
        RECT  1.9350 1.0450 2.0950 1.2850 ;
        RECT  1.1400 1.2750 2.0550 1.3950 ;
        RECT  1.1400 1.0550 1.2600 1.3950 ;
        RECT  0.7550 1.0550 1.2600 1.1750 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3550 1.2100 7.5950 1.3300 ;
        RECT  6.9950 1.2900 7.4750 1.4100 ;
        RECT  3.5500 1.5100 7.1150 1.6300 ;
        RECT  6.9950 1.2900 7.1150 1.6300 ;
        RECT  5.1400 1.2050 5.2600 1.6300 ;
        RECT  5.0200 1.2050 5.2600 1.3250 ;
        RECT  3.5500 1.2900 3.6700 1.6300 ;
        RECT  2.4900 1.2900 3.6700 1.4100 ;
        RECT  2.6350 1.2050 2.8750 1.4100 ;
        RECT  0.9000 1.5150 2.6100 1.6350 ;
        RECT  2.4900 1.2900 2.6100 1.6350 ;
        RECT  0.9000 1.2950 1.0200 1.6350 ;
        RECT  0.3900 1.2950 1.0200 1.4150 ;
        RECT  0.3900 0.8850 0.5100 1.4150 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.1940  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.9550 1.4700 9.0750 2.2100 ;
        RECT  8.7700 1.4650 9.0350 1.8750 ;
        RECT  8.9150 0.4850 9.0350 1.8750 ;
        RECT  1.4350 0.4850 9.0350 0.6050 ;
        RECT  0.5550 1.7550 9.0750 1.8750 ;
        RECT  8.1150 1.5000 8.2350 2.2100 ;
        RECT  7.2750 1.5300 7.3950 2.2100 ;
        RECT  6.4350 1.7500 6.5550 2.2100 ;
        RECT  5.5950 1.7500 5.7150 2.2100 ;
        RECT  4.7550 1.7500 4.8750 2.2100 ;
        RECT  3.9150 1.7500 4.0350 2.2100 ;
        RECT  3.0750 1.5300 3.1950 2.2100 ;
        RECT  2.2350 1.7550 2.3550 2.2100 ;
        RECT  1.3950 1.7550 1.5150 2.2100 ;
        RECT  0.5550 1.5350 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        RECT  7.6350 -0.1800 7.8750 0.3650 ;
        RECT  5.2500 -0.1800 5.4900 0.3650 ;
        RECT  2.4550 -0.1800 2.6950 0.3650 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        RECT  8.4750 1.9950 8.7150 2.1500 ;
        RECT  8.4750 1.9950 8.5950 2.7900 ;
        RECT  7.6350 1.9950 7.8750 2.1500 ;
        RECT  7.6350 1.9950 7.7550 2.7900 ;
        RECT  6.7950 1.9950 7.0350 2.1500 ;
        RECT  6.7950 1.9950 6.9150 2.7900 ;
        RECT  5.9550 1.9950 6.1950 2.1500 ;
        RECT  5.9550 1.9950 6.0750 2.7900 ;
        RECT  5.1150 1.9950 5.3550 2.1500 ;
        RECT  5.1150 1.9950 5.2350 2.7900 ;
        RECT  4.2750 1.9950 4.5150 2.1500 ;
        RECT  4.2750 1.9950 4.3950 2.7900 ;
        RECT  3.4350 1.9950 3.6750 2.1500 ;
        RECT  3.4350 1.9950 3.5550 2.7900 ;
        RECT  2.5950 1.9950 2.8350 2.1500 ;
        RECT  2.5950 1.9950 2.7150 2.7900 ;
        RECT  1.7550 1.9950 1.9950 2.1500 ;
        RECT  1.7550 1.9950 1.8750 2.7900 ;
        RECT  0.9150 1.9950 1.1550 2.1500 ;
        RECT  0.9150 1.9950 1.0350 2.7900 ;
        RECT  0.1350 1.4650 0.2550 2.7900 ;
        END
    END VDD
END NAND3X8

MACRO NAND3X6
    CLASS CORE ;
    FOREIGN NAND3X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9950 1.0550 6.2750 1.1750 ;
        RECT  5.9950 0.8200 6.1150 1.1750 ;
        RECT  4.1400 0.8200 6.1150 0.9400 ;
        RECT  3.9950 0.8400 4.2600 0.9600 ;
        RECT  3.3450 1.0350 4.1150 1.1550 ;
        RECT  3.9950 0.8400 4.1150 1.1550 ;
        RECT  3.5750 1.0350 3.8150 1.1750 ;
        RECT  3.3450 0.8200 3.4650 1.1550 ;
        RECT  2.0200 0.8200 3.4650 0.9400 ;
        RECT  1.7550 0.9400 2.1400 1.0900 ;
        RECT  1.5750 1.0550 1.8750 1.1750 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3950 1.0800 7.1950 1.2000 ;
        RECT  6.7400 0.8850 6.8900 1.2000 ;
        RECT  5.7550 1.2950 6.5150 1.4150 ;
        RECT  6.3950 1.0800 6.5150 1.4150 ;
        RECT  5.7550 1.0800 5.8750 1.4150 ;
        RECT  5.3000 1.0800 5.8750 1.2000 ;
        RECT  4.7000 1.0600 5.4200 1.1800 ;
        RECT  4.2350 1.0800 4.8200 1.2000 ;
        RECT  4.2350 1.0800 4.3550 1.3950 ;
        RECT  3.3350 1.2950 4.2500 1.4150 ;
        RECT  4.1300 1.2750 4.3550 1.3950 ;
        RECT  3.0700 1.2750 3.4550 1.3950 ;
        RECT  3.0700 1.0600 3.1900 1.3950 ;
        RECT  2.2750 1.0600 3.1900 1.1800 ;
        RECT  2.2750 1.0600 2.3950 1.3300 ;
        RECT  2.0100 1.2100 2.3950 1.3300 ;
        RECT  1.1400 1.2950 2.1300 1.4150 ;
        RECT  0.7550 1.2800 1.2600 1.4000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3700 1.1050 7.5550 1.3450 ;
        RECT  6.8600 1.3200 7.4900 1.4400 ;
        RECT  5.2700 1.5350 6.9800 1.6550 ;
        RECT  6.8600 1.3200 6.9800 1.6550 ;
        RECT  5.2700 1.3200 5.3900 1.6550 ;
        RECT  4.4750 1.3200 5.3900 1.4400 ;
        RECT  4.9400 1.3000 5.1800 1.4400 ;
        RECT  0.7100 1.5350 4.5950 1.6550 ;
        RECT  4.4750 1.3200 4.5950 1.6550 ;
        RECT  2.7100 1.3000 2.9500 1.6550 ;
        RECT  0.4450 1.5200 0.8300 1.6400 ;
        RECT  0.4450 1.2300 0.5650 1.6400 ;
        RECT  0.3250 1.2300 0.5650 1.4000 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.3781  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.7750 7.7950 1.8950 ;
        RECT  7.6750 0.5800 7.7950 1.8950 ;
        RECT  7.6100 1.4650 7.7950 1.8950 ;
        RECT  1.2950 0.5800 7.7950 0.7000 ;
        RECT  7.2750 1.5600 7.3950 2.2100 ;
        RECT  6.4350 1.7750 6.5550 2.2100 ;
        RECT  6.2350 0.4000 6.3550 0.9150 ;
        RECT  5.5950 1.7750 5.7150 2.2100 ;
        RECT  4.7550 1.5600 4.8750 2.2100 ;
        RECT  3.9150 1.7750 4.0350 2.2100 ;
        RECT  3.7550 0.4000 3.8750 0.9150 ;
        RECT  3.0750 1.7750 3.1950 2.2100 ;
        RECT  2.2350 1.7750 2.3550 2.2100 ;
        RECT  1.3950 1.7750 1.5150 2.2100 ;
        RECT  1.2950 0.4000 1.4150 0.9200 ;
        RECT  0.5550 1.7750 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  5.0750 0.3400 5.3150 0.4600 ;
        RECT  5.0750 -0.1800 5.1950 0.4600 ;
        RECT  2.5500 0.3400 2.7900 0.4600 ;
        RECT  2.5500 -0.1800 2.6700 0.4600 ;
        RECT  0.3350 -0.1800 0.4550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.6350 2.0150 7.8750 2.1500 ;
        RECT  7.6350 2.0150 7.7550 2.7900 ;
        RECT  6.7950 2.0150 7.0350 2.1500 ;
        RECT  6.7950 2.0150 6.9150 2.7900 ;
        RECT  5.9550 2.0150 6.1950 2.1500 ;
        RECT  5.9550 2.0150 6.0750 2.7900 ;
        RECT  5.1150 2.0150 5.3550 2.1500 ;
        RECT  5.1150 2.0150 5.2350 2.7900 ;
        RECT  4.2750 2.0150 4.5150 2.1500 ;
        RECT  4.2750 2.0150 4.3950 2.7900 ;
        RECT  3.4350 2.0150 3.6750 2.1500 ;
        RECT  3.4350 2.0150 3.5550 2.7900 ;
        RECT  2.5950 2.0150 2.8350 2.1500 ;
        RECT  2.5950 2.0150 2.7150 2.7900 ;
        RECT  1.7550 2.0150 1.9950 2.1500 ;
        RECT  1.7550 2.0150 1.8750 2.7900 ;
        RECT  0.9150 2.0150 1.1550 2.1500 ;
        RECT  0.9150 2.0150 1.0350 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
END NAND3X6

MACRO NAND3X4
    CLASS CORE ;
    FOREIGN NAND3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5750 0.9700 3.8150 1.0900 ;
        RECT  3.5750 0.8200 3.6950 1.0900 ;
        RECT  1.7550 0.8200 3.6950 0.9400 ;
        RECT  1.6150 0.9700 2.0150 1.0900 ;
        RECT  1.7550 0.8200 2.0150 1.0900 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4950 0.9600 4.6150 1.2000 ;
        RECT  4.4200 0.8850 4.5700 1.1450 ;
        RECT  3.9650 1.0250 4.6150 1.1450 ;
        RECT  3.3350 1.2100 4.0850 1.3300 ;
        RECT  3.9650 1.0250 4.0850 1.3300 ;
        RECT  3.0700 1.2000 3.4550 1.3200 ;
        RECT  3.0700 1.0600 3.1900 1.3200 ;
        RECT  2.2750 1.0600 3.1900 1.1800 ;
        RECT  1.2150 1.2100 2.3950 1.3300 ;
        RECT  2.2750 1.0600 2.3950 1.3300 ;
        RECT  1.2150 1.0800 1.3350 1.3300 ;
        RECT  0.7550 1.0800 1.3350 1.2000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7600 1.1050 4.9350 1.3450 ;
        RECT  4.4200 1.3200 4.8800 1.4400 ;
        RECT  0.9750 1.4500 4.5400 1.5700 ;
        RECT  4.4200 1.3200 4.5400 1.5700 ;
        RECT  2.7100 1.3000 2.9500 1.5700 ;
        RECT  0.9750 1.3200 1.0950 1.5700 ;
        RECT  0.4450 1.3200 1.0950 1.4400 ;
        RECT  0.3050 1.3000 0.6350 1.3800 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        RECT  0.3950 1.3200 1.0950 1.4200 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5232  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.6900 5.1750 1.8100 ;
        RECT  5.0550 0.5800 5.1750 1.8100 ;
        RECT  5.0000 1.4650 5.1750 1.8100 ;
        RECT  1.5350 0.5800 5.1750 0.7000 ;
        RECT  4.7550 1.5600 4.8750 2.2100 ;
        RECT  3.9150 1.6900 4.0350 2.2100 ;
        RECT  3.0750 1.6900 3.1950 2.2100 ;
        RECT  2.2350 1.6900 2.3550 2.2100 ;
        RECT  1.3950 1.6900 1.5150 2.2100 ;
        RECT  0.5550 1.5600 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.9750 0.3400 5.2150 0.4600 ;
        RECT  4.9750 -0.1800 5.0950 0.4600 ;
        RECT  2.5550 0.3400 2.7950 0.4600 ;
        RECT  2.5550 -0.1800 2.6750 0.4600 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  5.1750 1.9300 5.2950 2.7900 ;
        RECT  4.3350 1.9300 4.4550 2.7900 ;
        RECT  3.4950 1.9300 3.6150 2.7900 ;
        RECT  2.6550 1.9300 2.7750 2.7900 ;
        RECT  1.8150 1.9300 1.9350 2.7900 ;
        RECT  0.9750 1.9300 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
END NAND3X4

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2950 0.7500 2.4150 1.1700 ;
        RECT  0.3900 0.7500 2.4150 0.8700 ;
        RECT  0.4950 0.7500 0.6150 1.1700 ;
        RECT  0.3600 0.8850 0.6150 1.1450 ;
        RECT  0.3900 0.7500 0.6150 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.9900 2.0950 1.2300 ;
        RECT  1.8100 0.9900 1.9600 1.4350 ;
        RECT  0.7550 0.9900 2.0950 1.1100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2300 1.5550 1.4200 ;
        RECT  1.1750 1.2300 1.4350 1.4450 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7616  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5650 2.6550 1.6850 ;
        RECT  2.5350 0.5100 2.6550 1.6850 ;
        RECT  2.3350 1.5200 2.6550 1.6850 ;
        RECT  1.4350 0.5100 2.6550 0.6300 ;
        RECT  2.2350 1.5600 2.3550 2.2100 ;
        RECT  1.3950 1.5650 1.5150 2.2100 ;
        RECT  0.5550 1.5600 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.4550 -0.1800 2.6950 0.3900 ;
        RECT  0.2750 0.4600 0.5150 0.5800 ;
        RECT  0.2750 -0.1800 0.3950 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.6550 1.8050 2.7750 2.7900 ;
        RECT  1.8150 1.8050 1.9350 2.7900 ;
        RECT  0.9750 1.8050 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
END NAND3X2

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.8250 0.8200 1.2400 ;
        RECT  0.6500 0.5950 0.8000 0.9950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7600 0.5100 1.2150 ;
        RECT  0.3800 0.7600 0.5000 1.2400 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 0.8850 1.1750 1.2050 ;
        RECT  0.9400 0.8850 1.0900 1.2100 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5104  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.3600 1.5150 2.2100 ;
        RECT  1.2950 0.6450 1.4150 1.7250 ;
        RECT  1.1950 0.5250 1.3150 0.7650 ;
        RECT  1.2300 1.3600 1.5150 1.7250 ;
        RECT  0.5550 1.3600 1.5150 1.4800 ;
        RECT  0.5550 1.3600 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.2200 -0.1800 0.3400 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.6000 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
END NAND3X1

MACRO NAND3BXL
    CLASS CORE ;
    FOREIGN NAND3BXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0400 0.5100 1.5100 ;
        RECT  0.3600 1.0400 0.4800 1.5400 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8100 1.0200 0.9350 1.2600 ;
        RECT  0.6500 1.0200 0.9350 1.1450 ;
        RECT  0.6500 0.8850 0.8050 1.1450 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5150 1.3550 1.6700 1.7350 ;
        RECT  1.4800 1.3550 1.6700 1.7250 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9150 1.8400 1.1550 1.9600 ;
        RECT  0.9150 1.6600 1.0350 1.9600 ;
        RECT  0.1200 1.6600 1.0350 1.7800 ;
        RECT  0.1200 0.8000 0.4550 0.9200 ;
        RECT  0.3350 0.6800 0.4550 0.9200 ;
        RECT  0.1350 1.6600 0.2550 2.0200 ;
        RECT  0.0700 1.4650 0.2400 1.7250 ;
        RECT  0.1200 0.8000 0.2400 1.7800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.2950 -0.1800 1.4150 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.3950 1.9000 1.5150 2.7900 ;
        RECT  0.5550 1.9000 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 2.0200 1.8150 2.0200 1.8150 1.9000 1.7900 1.9000 1.7900 1.2350 1.1500 1.2350
                 1.1500 1.1150 1.7150 1.1150 1.7150 0.6800 1.8350 0.6800 1.8350 0.9950 1.9100 0.9950
                 1.9100 1.7800 1.9350 1.7800 ;
    END
END NAND3BXL

MACRO NAND3BX4
    CLASS CORE ;
    FOREIGN NAND3BX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5750 0.9700 3.8150 1.0900 ;
        RECT  3.5750 0.8200 3.6950 1.0900 ;
        RECT  2.2000 0.8200 3.6950 0.9400 ;
        RECT  1.6150 0.9700 2.3200 1.0900 ;
        RECT  2.2000 0.8200 2.3200 1.0900 ;
        RECT  1.7550 0.9400 2.0150 1.0900 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0850 0.9850 5.4150 1.1200 ;
        RECT  4.9450 0.9400 5.2050 1.1050 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9350 1.0800 4.6750 1.2000 ;
        RECT  3.2350 1.2100 4.0550 1.3300 ;
        RECT  3.9350 1.0800 4.0550 1.3300 ;
        RECT  3.2350 1.0600 3.3550 1.3300 ;
        RECT  2.4400 1.0600 3.3550 1.1800 ;
        RECT  1.1150 1.2100 2.5600 1.3300 ;
        RECT  2.4400 1.0600 2.5600 1.3300 ;
        RECT  1.1150 1.0800 1.2350 1.3300 ;
        RECT  0.8850 0.9400 1.1450 1.2000 ;
        RECT  0.7550 1.0800 1.2350 1.2000 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5232  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7550 1.5600 4.8750 2.2100 ;
        RECT  0.2550 1.6900 4.8750 1.8100 ;
        RECT  3.9150 1.6900 4.0350 2.2100 ;
        RECT  0.2550 0.5800 3.8950 0.7000 ;
        RECT  3.0750 1.6900 3.1950 2.2100 ;
        RECT  2.2350 1.6900 2.3550 2.2100 ;
        RECT  1.3950 1.6900 1.5150 2.2100 ;
        RECT  0.5550 1.5600 0.6750 2.2100 ;
        RECT  0.0700 1.4650 0.3750 1.7250 ;
        RECT  0.2550 0.5800 0.3750 1.8100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  4.9750 -0.1800 5.0950 0.6400 ;
        RECT  2.4950 0.3400 2.7350 0.4600 ;
        RECT  2.4950 -0.1800 2.6150 0.4600 ;
        RECT  0.2150 0.3400 0.4550 0.4600 ;
        RECT  0.2150 -0.1800 0.3350 0.4600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1750 1.5600 5.2950 2.7900 ;
        RECT  4.3350 1.9300 4.4550 2.7900 ;
        RECT  3.4950 1.9300 3.6150 2.7900 ;
        RECT  2.6550 1.9300 2.7750 2.7900 ;
        RECT  1.8150 1.9300 1.9350 2.7900 ;
        RECT  0.9750 1.9300 1.0950 2.7900 ;
        RECT  0.1350 1.9300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7150 2.2100 5.5950 2.2100 5.5950 1.5200 5.5350 1.5200 5.5350 1.4000 4.9150 1.4000
                 4.9150 1.4400 4.3850 1.4400 4.3850 1.5700 0.8200 1.5700 0.8200 1.4400 0.4950 1.4400
                 0.4950 1.2000 0.6150 1.2000 0.6150 1.3200 0.9400 1.3200 0.9400 1.4500 2.8350 1.4500
                 2.8350 1.3000 3.0750 1.3000 3.0750 1.4500 4.2650 1.4500 4.2650 1.3200 4.7950 1.3200
                 4.7950 1.2800 5.5350 1.2800 5.5350 0.8650 5.3950 0.8650 5.3950 0.5900 5.5150 0.5900
                 5.5150 0.7450 5.6550 0.7450 5.6550 1.4000 5.7150 1.4000 ;
    END
END NAND3BX4

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7650 0.9900 2.8850 1.4200 ;
        RECT  2.6800 1.0250 2.8300 1.4400 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  2.0250 0.9900 2.2200 1.2300 ;
        RECT  0.8050 0.9900 2.2200 1.1100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2300 1.4350 1.5000 ;
        RECT  1.1250 1.2300 1.4350 1.4800 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7616  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2850 1.5600 2.4050 2.2100 ;
        RECT  0.3050 1.6200 2.4050 1.7400 ;
        RECT  1.4450 1.6200 1.5650 2.2100 ;
        RECT  0.3050 0.5100 1.5250 0.6300 ;
        RECT  0.6050 1.5600 0.7250 2.2100 ;
        RECT  0.3050 1.5600 0.7250 1.7400 ;
        RECT  0.3050 1.5200 0.5650 1.7400 ;
        RECT  0.3050 0.5100 0.4250 1.7400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.4450 0.4600 2.6850 0.5800 ;
        RECT  2.4450 -0.1800 2.5650 0.5800 ;
        RECT  0.2650 -0.1800 0.5050 0.3900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.7050 1.5600 2.8250 2.7900 ;
        RECT  1.8650 1.8600 1.9850 2.7900 ;
        RECT  1.0250 1.8600 1.1450 2.7900 ;
        RECT  0.1850 1.8600 0.3050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.3050 1.8000 3.1850 1.8000 3.1850 1.6800 3.0050 1.6800 3.0050 0.8700 2.5600 0.8700
                 2.5600 1.1700 2.4400 1.1700 2.4400 0.8700 0.6650 0.8700 0.6650 1.1700 0.5450 1.1700
                 0.5450 0.7500 2.9850 0.7500 2.9850 0.5900 3.1050 0.5900 3.1050 0.7100 3.1250 0.7100
                 3.1250 1.5600 3.3050 1.5600 ;
    END
END NAND3BX2

MACRO NAND3BX1
    CLASS CORE ;
    FOREIGN NAND3BX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7850 0.5100 1.2400 ;
        RECT  0.3600 0.7600 0.4800 1.2400 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8150 0.9300 0.9350 1.1700 ;
        RECT  0.6500 0.9300 0.9350 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.0000 1.6700 1.5000 ;
        RECT  1.5200 1.0000 1.6700 1.4700 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5104  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9750 1.3600 1.0950 2.2100 ;
        RECT  0.1200 1.3600 1.0950 1.4800 ;
        RECT  0.1200 0.5200 0.4550 0.6400 ;
        RECT  0.3350 0.4000 0.4550 0.6400 ;
        RECT  0.1350 1.3600 0.2550 2.2100 ;
        RECT  0.0700 1.1750 0.2400 1.4350 ;
        RECT  0.1200 0.5200 0.2400 1.4800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.2950 -0.1800 1.4150 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.3950 1.6200 1.5150 2.7900 ;
        RECT  0.5550 1.6000 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9950 1.8000 1.8750 1.8000 1.8750 1.6800 1.7900 1.6800 1.7900 0.8800 1.4000 0.8800
                 1.4000 1.1100 1.1500 1.1100 1.1500 0.9900 1.2800 0.9900 1.2800 0.7600 1.7750 0.7600
                 1.7750 0.5900 1.8950 0.5900 1.8950 0.7100 1.9100 0.7100 1.9100 1.5600 1.9950 1.5600 ;
    END
END NAND3BX1

MACRO NAND2XL
    CLASS CORE ;
    FOREIGN NAND2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.1600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5850 1.1750 0.8000 1.4350 ;
        RECT  0.6100 1.0550 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.3600 1.4400 ;
        RECT  0.2400 1.0400 0.3600 1.4400 ;
        RECT  0.0700 1.1750 0.2200 1.5650 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4800 1.5550 1.0400 1.6750 ;
        RECT  0.9200 0.8000 1.0400 1.6750 ;
        RECT  0.6500 0.6800 0.9400 0.8550 ;
        RECT  0.6800 0.8000 1.0400 0.9200 ;
        RECT  0.6500 0.5950 0.8000 0.8550 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.1600 0.1800 ;
        RECT  0.1800 -0.1800 0.3000 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.1600 2.7900 ;
        RECT  0.9050 2.0200 1.0250 2.7900 ;
        RECT  0.1350 2.0200 0.2550 2.7900 ;
        END
    END VDD
END NAND2XL

MACRO NAND2X8
    CLASS CORE ;
    FOREIGN NAND2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8550 1.0500 5.0950 1.1700 ;
        RECT  0.3050 0.9650 4.9750 1.0850 ;
        RECT  3.6950 0.9650 3.9350 1.1700 ;
        RECT  1.8150 0.9650 2.0550 1.1700 ;
        RECT  0.4350 0.9650 0.6750 1.1750 ;
        RECT  0.3050 0.9400 0.5650 1.0900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3750 1.1900 5.8350 1.3100 ;
        RECT  1.1750 1.2900 5.4950 1.4100 ;
        RECT  5.2350 1.2300 5.8350 1.3100 ;
        RECT  4.0550 1.2100 4.2950 1.4100 ;
        RECT  2.8750 1.2050 3.1150 1.4100 ;
        RECT  1.0550 1.2050 1.2950 1.3250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.2732  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5300 6.0750 1.6500 ;
        RECT  5.9550 0.7100 6.0750 1.6500 ;
        RECT  5.8700 1.4650 6.0200 1.7250 ;
        RECT  0.9150 0.7100 6.0750 0.8300 ;
        RECT  5.5950 1.5300 5.7150 2.2100 ;
        RECT  4.7550 1.5300 4.8750 2.2100 ;
        RECT  3.9150 1.5300 4.0350 2.2100 ;
        RECT  3.0750 1.5300 3.1950 2.2100 ;
        RECT  2.2350 1.5300 2.3550 2.2100 ;
        RECT  1.3950 1.5300 1.5150 2.2100 ;
        RECT  0.5550 1.4650 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.1150 0.4600 5.3550 0.5800 ;
        RECT  5.1150 -0.1800 5.2350 0.5800 ;
        RECT  3.5550 0.4600 3.7950 0.5800 ;
        RECT  3.5550 -0.1800 3.6750 0.5800 ;
        RECT  1.5550 0.4600 1.7950 0.5800 ;
        RECT  1.5550 -0.1800 1.6750 0.5800 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  6.0150 1.8450 6.1350 2.7900 ;
        RECT  5.1750 1.7700 5.2950 2.7900 ;
        RECT  4.3350 1.7700 4.4550 2.7900 ;
        RECT  3.4950 1.7700 3.6150 2.7900 ;
        RECT  2.6550 1.7700 2.7750 2.7900 ;
        RECT  1.8150 1.7700 1.9350 2.7900 ;
        RECT  0.9750 1.7700 1.0950 2.7900 ;
        RECT  0.1350 1.4650 0.2550 2.7900 ;
        END
    END VDD
END NAND2X8

MACRO NAND2X6
    CLASS CORE ;
    FOREIGN NAND2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9150 0.9900 5.0350 1.3450 ;
        RECT  0.6500 0.9900 5.0350 1.1100 ;
        RECT  3.4250 0.9900 3.6650 1.1950 ;
        RECT  1.9150 0.9900 2.1550 1.1950 ;
        RECT  0.4350 1.0800 0.8000 1.2000 ;
        RECT  0.6500 0.8850 0.8000 1.2000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.3000 4.1750 1.4200 ;
        RECT  3.7850 1.2300 4.0450 1.4200 ;
        RECT  1.2950 1.3150 3.9050 1.4350 ;
        RECT  2.6550 1.3000 2.8950 1.4350 ;
        RECT  1.1750 1.2800 1.4150 1.4000 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.7541  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5550 5.2750 1.6750 ;
        RECT  5.1550 0.7500 5.2750 1.6750 ;
        RECT  5.0000 1.4650 5.2750 1.6750 ;
        RECT  0.9750 0.7500 5.2750 0.8700 ;
        RECT  5.0000 1.4650 5.1500 1.7250 ;
        RECT  4.7550 1.5550 4.8750 2.2100 ;
        RECT  4.1350 0.4000 4.2550 0.8700 ;
        RECT  3.9150 1.5550 4.0350 2.2100 ;
        RECT  3.0750 1.5550 3.1950 2.2100 ;
        RECT  2.8550 0.4000 2.9750 0.8700 ;
        RECT  2.2350 1.5550 2.3550 2.2100 ;
        RECT  1.3950 1.5550 1.5150 2.2100 ;
        RECT  0.9750 0.4000 1.0950 0.8700 ;
        RECT  0.5550 1.5550 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  3.4350 0.4600 3.6750 0.6300 ;
        RECT  3.4350 -0.1800 3.5550 0.6300 ;
        RECT  1.6550 0.4600 1.8950 0.6300 ;
        RECT  1.6550 -0.1800 1.7750 0.6300 ;
        RECT  0.3350 -0.1800 0.4550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  5.1750 1.8450 5.2950 2.7900 ;
        RECT  4.3350 1.7950 4.4550 2.7900 ;
        RECT  3.4950 1.7950 3.6150 2.7900 ;
        RECT  2.6550 1.7950 2.7750 2.7900 ;
        RECT  1.8150 1.7950 1.9350 2.7900 ;
        RECT  0.9750 1.7950 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
END NAND2X6

MACRO NAND2X4
    CLASS CORE ;
    FOREIGN NAND2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4350 0.9900 3.3150 1.1100 ;
        RECT  0.5950 0.9400 0.8550 1.1100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.2300 2.5950 1.3800 ;
        RECT  1.1750 1.2300 2.5950 1.3500 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1072  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5000 3.5550 1.6200 ;
        RECT  3.4350 0.7000 3.5550 1.6200 ;
        RECT  3.2050 1.2300 3.5550 1.3800 ;
        RECT  1.3350 0.7000 3.5550 0.8200 ;
        RECT  3.0750 1.5000 3.1950 2.2100 ;
        RECT  2.4950 0.6500 2.7350 0.8200 ;
        RECT  2.2350 1.5000 2.3550 2.2100 ;
        RECT  1.3950 1.5000 1.5150 2.2100 ;
        RECT  1.2150 0.6500 1.4550 0.7700 ;
        RECT  0.5550 1.5000 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.1350 0.4600 3.3750 0.5800 ;
        RECT  3.1350 -0.1800 3.2550 0.5800 ;
        RECT  1.8550 0.4600 2.0950 0.5800 ;
        RECT  1.8550 -0.1800 1.9750 0.5800 ;
        RECT  0.6350 -0.1800 0.7550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.4950 1.7400 3.6150 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
END NAND2X4

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5350 0.9900 1.7750 1.1100 ;
        RECT  0.5950 0.9400 1.6550 0.9900 ;
        RECT  0.7350 0.8700 1.6550 0.9900 ;
        RECT  0.5750 0.9900 0.8550 1.1100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.1100 1.3800 1.5800 ;
        RECT  1.2300 1.1100 1.3500 1.6100 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5536  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6950 1.7300 2.0150 1.8500 ;
        RECT  1.8950 0.6300 2.0150 1.8500 ;
        RECT  1.7550 1.2300 2.0150 1.3800 ;
        RECT  1.0550 0.6300 2.0150 0.7500 ;
        RECT  1.5350 1.5600 1.6550 2.2100 ;
        RECT  0.6950 1.5600 0.8150 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.7550 0.3900 1.9950 0.5100 ;
        RECT  1.7550 -0.1800 1.8750 0.5100 ;
        RECT  0.4750 -0.1800 0.5950 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.9550 1.9700 2.0750 2.7900 ;
        RECT  1.1150 1.9700 1.2350 2.7900 ;
        RECT  0.2750 1.5600 0.3950 2.7900 ;
        END
    END VDD
END NAND2X2

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.4500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 0.5950 0.8000 1.2000 ;
        RECT  0.6500 0.5950 0.8000 1.0200 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.8250 0.5100 1.2000 ;
        RECT  0.3600 0.8250 0.4800 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3284  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9200 1.1750 1.0900 1.4350 ;
        RECT  0.6200 1.3200 1.0400 1.4400 ;
        RECT  0.9200 0.6200 1.0400 1.4400 ;
        RECT  0.6200 1.3200 0.7400 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.4500 0.1800 ;
        RECT  0.2000 -0.1800 0.3200 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.4500 2.7900 ;
        RECT  1.0400 1.5600 1.1600 2.7900 ;
        RECT  0.2000 1.5600 0.3200 2.7900 ;
        END
    END VDD
END NAND2X1

MACRO NAND2BXL
    CLASS CORE ;
    FOREIGN NAND2BXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4900 0.8650 0.6350 1.1050 ;
        RECT  0.3600 0.8850 0.5350 1.1450 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.2750 1.3650 ;
        RECT  1.1550 1.1250 1.2750 1.3650 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.3150 0.6750 1.6850 ;
        RECT  0.0700 1.3150 0.6750 1.4350 ;
        RECT  0.1200 0.6450 0.3700 0.7650 ;
        RECT  0.2500 0.5250 0.3700 0.7650 ;
        RECT  0.0700 1.1750 0.2400 1.4350 ;
        RECT  0.1200 0.6450 0.2400 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9700 -0.1800 1.0900 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.0050 2.0850 1.1250 2.7900 ;
        RECT  0.1350 1.5650 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6050 1.6850 1.4850 1.6850 1.4850 1.5650 1.3950 1.5650 1.3950 1.0050 1.0350 1.0050
                 1.0350 1.0450 0.7550 1.0450 0.7550 0.9250 0.9150 0.9250 0.9150 0.8850 1.3950 0.8850
                 1.3950 0.7650 1.3900 0.7650 1.3900 0.5250 1.5100 0.5250 1.5100 0.6450 1.5150 0.6450
                 1.5150 1.4450 1.6050 1.4450 ;
    END
END NAND2BXL

MACRO NAND2BX4
    CLASS CORE ;
    FOREIGN NAND2BX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 1.3300 3.7000 1.7250 ;
        RECT  3.5800 1.2400 3.7000 1.7250 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.2600 2.7800 1.3800 ;
        RECT  2.3350 1.2300 2.5950 1.3800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1072  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0800 1.5000 3.2000 2.2100 ;
        RECT  0.2000 1.5000 3.2000 1.6200 ;
        RECT  2.7000 0.6500 2.9400 0.7700 ;
        RECT  0.2000 0.7000 2.8200 0.8200 ;
        RECT  2.2400 1.5000 2.3600 2.2100 ;
        RECT  1.4200 0.6500 1.6600 0.8200 ;
        RECT  1.4000 1.5000 1.5200 2.2100 ;
        RECT  0.5600 1.5000 0.6800 2.2100 ;
        RECT  0.2000 1.2300 0.5650 1.3800 ;
        RECT  0.2000 0.7000 0.3200 1.6200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.4000 -0.1800 3.5200 0.6400 ;
        RECT  2.0600 0.4600 2.3000 0.5800 ;
        RECT  2.0600 -0.1800 2.1800 0.5800 ;
        RECT  0.7800 0.4600 1.0200 0.5800 ;
        RECT  0.7800 -0.1800 0.9000 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.5000 1.8450 3.6200 2.7900 ;
        RECT  2.6600 1.7400 2.7800 2.7900 ;
        RECT  1.8200 1.7400 1.9400 2.7900 ;
        RECT  0.9800 1.7400 1.1000 2.7900 ;
        RECT  0.1400 1.7400 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.0400 2.2100 3.9200 2.2100 3.9200 1.6800 3.8200 1.6800 3.8200 1.1100 0.4400 1.1100
                 0.4400 0.9900 3.8200 0.9900 3.8200 0.5900 3.9400 0.5900 3.9400 1.5600 4.0400 1.5600 ;
    END
END NAND2BX4

MACRO NAND2BX2
    CLASS CORE ;
    FOREIGN NAND2BX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2050 1.2650 1.3950 ;
        RECT  0.8850 1.1800 1.1450 1.3950 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0150 1.2400 2.1350 1.4800 ;
        RECT  1.8400 1.3600 2.1350 1.4800 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5536  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.5150 1.5150 2.2100 ;
        RECT  0.1950 1.5150 1.5150 1.6350 ;
        RECT  1.1150 0.6500 1.3550 0.7700 ;
        RECT  0.1950 0.7000 1.2350 0.8200 ;
        RECT  0.5550 1.5150 0.6750 2.2100 ;
        RECT  0.1950 0.7000 0.3150 1.6350 ;
        RECT  0.0700 0.8850 0.3150 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8150 -0.1800 1.9350 0.6400 ;
        RECT  0.4750 0.4600 0.7150 0.5800 ;
        RECT  0.4750 -0.1800 0.5950 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8150 1.8450 1.9350 2.7900 ;
        RECT  0.9750 1.7550 1.0950 2.7900 ;
        RECT  0.1350 1.7550 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4150 1.8000 2.2950 1.8000 2.2950 1.0600 1.8350 1.0600 1.8350 1.1100 1.5950 1.1100
                 1.5950 1.0600 0.7650 1.0600 0.7650 1.1100 0.4350 1.1100 0.4350 0.9900 0.6450 0.9900
                 0.6450 0.9400 2.2950 0.9400 2.2950 0.5900 2.4150 0.5900 ;
    END
END NAND2BX2

MACRO NAND2BX1
    CLASS CORE ;
    FOREIGN NAND2BX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.7600 0.5100 1.2400 ;
        RECT  0.3600 0.7600 0.5100 1.2150 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.0000 1.3800 1.5000 ;
        RECT  1.2300 1.0000 1.3800 1.4700 ;
        END
    END AN
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3284  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6200 1.3600 0.7400 2.2100 ;
        RECT  0.1200 1.3600 0.7400 1.4800 ;
        RECT  0.1200 0.5200 0.4600 0.6400 ;
        RECT  0.3400 0.4000 0.4600 0.6400 ;
        RECT  0.0700 1.1750 0.2400 1.4350 ;
        RECT  0.1200 0.5200 0.2400 1.4800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9800 -0.1800 1.1000 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.0400 1.6200 1.1600 2.7900 ;
        RECT  0.2000 1.6000 0.3200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6200 1.7400 1.5800 1.7400 1.5800 1.8600 1.4600 1.8600 1.4600 1.6200 1.5000 1.6200
                 1.5000 0.8800 1.1100 0.8800 1.1100 1.0900 0.8400 1.0900 0.8400 0.9700 0.9900 0.9700
                 0.9900 0.7600 1.4600 0.7600 1.4600 0.5900 1.5800 0.5900 1.5800 0.7100 1.6200 0.7100 ;
    END
END NAND2BX1

MACRO MXI4XL
    CLASS CORE ;
    FOREIGN MXI4XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 0.4800 2.4550 1.0800 ;
        RECT  2.3150 0.9600 2.4350 1.4700 ;
        RECT  0.6800 0.4800 2.4550 0.6000 ;
        RECT  1.8350 0.4000 2.0750 0.6000 ;
        RECT  0.6800 1.0000 0.8400 1.2400 ;
        RECT  0.6800 0.4800 0.8000 1.2400 ;
        RECT  0.6500 0.5950 0.8000 0.8550 ;
        END
    END S1
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0350 1.2600 3.2750 1.4600 ;
        RECT  2.9150 1.1550 3.1750 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0750 1.5100 4.5350 1.6500 ;
        RECT  4.0750 1.5000 4.3350 1.6700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6550 1.4400 4.9150 1.6700 ;
        RECT  4.6950 1.2600 4.8150 1.6700 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9550 1.5500 6.2350 1.7000 ;
        RECT  5.8150 1.5000 6.0750 1.6850 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.1752  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.9733  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7750 1.2600 6.5750 1.3800 ;
        RECT  6.1050 1.2300 6.3650 1.3800 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6600 0.2550 1.5800 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  6.2350 -0.1800 6.3550 0.3800 ;
        RECT  4.5550 -0.1800 4.6750 0.3800 ;
        RECT  2.8550 -0.1800 2.9750 0.8600 ;
        RECT  1.3100 -0.1800 1.5500 0.3200 ;
        RECT  0.5550 -0.1800 0.7950 0.3200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  6.1350 1.9600 6.2550 2.7900 ;
        RECT  4.6850 2.0300 4.8050 2.7900 ;
        RECT  4.5650 2.0300 4.8050 2.1500 ;
        RECT  2.8950 2.1400 3.0150 2.7900 ;
        RECT  1.2550 1.9100 1.3750 2.7900 ;
        RECT  1.1350 1.9100 1.3750 2.0300 ;
        RECT  0.5550 2.0400 0.7950 2.1600 ;
        RECT  0.5550 2.0400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.8250 0.9000 6.8150 0.9000 6.8150 1.6200 6.6750 1.6200 6.6750 2.0800 6.5550 2.0800
                 6.5550 1.5000 6.6950 1.5000 6.6950 0.7800 6.7050 0.7800 6.7050 0.6200 5.9950 0.6200
                 5.9950 0.5400 5.4150 0.5400 5.4150 1.6700 5.2950 1.6700 5.2950 0.6200 4.3100 0.6200
                 4.3100 0.5600 3.6350 0.5600 3.6350 1.5400 3.3950 1.5400 3.3950 1.4200 3.5150 1.4200
                 3.5150 0.4400 3.9350 0.4400 3.9350 0.3600 4.1750 0.3600 4.1750 0.4400 4.4300 0.4400
                 4.4300 0.5000 5.2950 0.5000 5.2950 0.4200 5.6150 0.4200 5.6150 0.4000 5.8550 0.4000
                 5.8550 0.4200 6.1150 0.4200 6.1150 0.5000 6.8250 0.5000 ;
        POLYGON  5.6550 1.9600 5.5750 1.9600 5.5750 2.0800 5.4550 2.0800 5.4550 1.9600 4.9250 1.9600
                 4.9250 1.9100 4.2500 1.9100 4.2500 2.2500 3.3350 2.2500 3.3350 2.1300 3.1350 2.1300
                 3.1350 2.0200 2.6750 2.0200 2.6750 2.2500 2.5550 2.2500 2.5550 1.9000 3.2550 1.9000
                 3.2550 2.0100 3.4550 2.0100 3.4550 2.1300 4.1300 2.1300 4.1300 1.7900 5.0450 1.7900
                 5.0450 1.8400 5.5350 1.8400 5.5350 0.6600 5.6550 0.6600 ;
        POLYGON  5.1750 1.1600 4.9350 1.1600 4.9350 1.1400 4.1150 1.1400 4.1150 1.3800 3.9950 1.3800
                 3.9950 1.0200 5.1750 1.0200 ;
        POLYGON  4.0350 0.8000 3.8750 0.8000 3.8750 1.8900 3.7150 1.8900 3.7150 2.0100 3.5950 2.0100
                 3.5950 1.8900 3.3750 1.8900 3.3750 1.7800 2.4350 1.7800 2.4350 2.1100 1.7350 2.1100
                 1.7350 2.2500 1.4950 2.2500 1.4950 2.1300 1.6150 2.1300 1.6150 1.9900 2.3150 1.9900
                 2.3150 1.6600 3.4950 1.6600 3.4950 1.7700 3.7550 1.7700 3.7550 0.6800 4.0350 0.6800 ;
        POLYGON  2.2150 0.8400 2.1950 0.8400 2.1950 1.7500 2.1750 1.7500 2.1750 1.8700 2.0550 1.8700
                 2.0550 1.7600 0.3800 1.7600 0.3800 1.0200 0.5000 1.0200 0.5000 1.6400 2.0550 1.6400
                 2.0550 1.6300 2.0750 1.6300 2.0750 0.8400 1.9750 0.8400 1.9750 0.7200 2.2150 0.7200 ;
        POLYGON  1.9550 1.4700 1.2250 1.4700 1.2250 1.5200 0.9850 1.5200 0.9850 1.4000 1.0400 1.4000
                 1.0400 0.8400 0.9200 0.8400 0.9200 0.7200 1.1600 0.7200 1.1600 1.3500 1.8350 1.3500
                 1.8350 1.2300 1.9550 1.2300 ;
    END
END MXI4XL

MACRO MXI4X4
    CLASS CORE ;
    FOREIGN MXI4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.2904  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.6133  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0350 1.2000 1.1550 1.4400 ;
        RECT  0.3900 1.2000 1.1550 1.3200 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        RECT  0.3900 1.2000 0.5100 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.4400 0.8350 1.8500 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1150 1.2900 2.2550 1.6850 ;
        RECT  2.0800 1.3400 2.2500 1.7250 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.3100 2.6150 1.7250 ;
        RECT  2.4950 1.2900 2.6150 1.7250 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8400 1.3600 4.0050 1.7250 ;
        RECT  3.8350 1.2800 3.9700 1.6500 ;
        END
    END D
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6952  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7150 1.5700 7.9550 1.6900 ;
        RECT  6.7550 0.9500 7.9550 1.0700 ;
        RECT  7.8350 0.6000 7.9550 1.0700 ;
        RECT  7.7150 0.9500 7.8350 1.6900 ;
        RECT  7.6100 0.9500 7.8350 1.4350 ;
        RECT  6.7550 1.5700 6.9950 1.6900 ;
        RECT  6.8550 0.9500 6.9750 1.6900 ;
        RECT  6.7550 0.6000 6.8750 1.0700 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1350 1.5200 8.6550 1.6400 ;
        RECT  7.4800 1.8100 8.3950 1.9300 ;
        RECT  8.2750 1.5200 8.3950 1.9300 ;
        RECT  8.1350 1.5200 8.3950 1.6700 ;
        RECT  7.4800 1.8100 7.6000 2.1700 ;
        RECT  5.8900 2.0500 7.6000 2.1700 ;
        RECT  4.5750 2.1300 6.0100 2.2500 ;
        RECT  4.5750 1.3300 4.6950 2.2500 ;
        END
    END S1
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.3150 -0.1800 8.4350 0.8400 ;
        RECT  7.2350 0.4700 7.4750 0.5900 ;
        RECT  7.3550 -0.1800 7.4750 0.5900 ;
        RECT  6.2750 -0.1800 6.3950 0.7900 ;
        RECT  4.0850 -0.1800 4.2050 0.9200 ;
        RECT  2.3550 -0.1800 2.4750 0.3800 ;
        RECT  0.4950 0.7200 0.7350 0.8400 ;
        RECT  0.4950 -0.1800 0.6150 0.8400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.1950 2.0500 8.4350 2.1700 ;
        RECT  8.1950 2.0500 8.3150 2.7900 ;
        RECT  7.2350 2.2900 7.4750 2.7900 ;
        RECT  6.1300 2.2900 6.3700 2.7900 ;
        RECT  3.7000 2.0850 3.9400 2.2050 ;
        RECT  3.7000 2.0850 3.8200 2.7900 ;
        RECT  2.0550 2.0850 2.2950 2.2050 ;
        RECT  2.0550 2.0850 2.1750 2.7900 ;
        RECT  0.7150 1.9700 0.8350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.8950 1.8800 8.8550 1.8800 8.8550 2.0400 8.7350 2.0400 8.7350 1.7600 8.7750 1.7600
                 8.7750 1.0800 8.0750 1.0800 8.0750 0.4800 7.7150 0.4800 7.7150 0.8300 6.9950 0.8300
                 6.9950 0.4800 6.6350 0.4800 6.6350 1.6900 5.4350 1.6900 5.4350 1.5400 4.8950 1.5400
                 4.8950 1.0200 5.0150 1.0200 5.0150 1.4200 5.4350 1.4200 5.4350 1.3000 5.5550 1.3000
                 5.5550 1.5700 6.5150 1.5700 6.5150 0.3600 7.1150 0.3600 7.1150 0.7100 7.5950 0.7100
                 7.5950 0.3600 8.1950 0.3600 8.1950 0.9600 8.6050 0.9600 8.6050 0.7200 8.7350 0.7200
                 8.7350 0.6000 8.8550 0.6000 8.8550 0.7200 8.8950 0.7200 ;
        POLYGON  7.2350 1.9300 5.3150 1.9300 5.3150 2.0100 5.1950 2.0100 5.1950 1.6700 5.3150 1.6700
                 5.3150 1.8100 7.1150 1.8100 7.1150 1.4300 7.0950 1.4300 7.0950 1.1900 7.2150 1.1900
                 7.2150 1.3100 7.2350 1.3100 ;
        POLYGON  6.3950 1.4500 5.6750 1.4500 5.6750 1.0100 5.1350 1.0100 5.1350 0.8900 4.9550 0.8900
                 4.9550 0.6500 5.0750 0.6500 5.0750 0.7700 5.2550 0.7700 5.2550 0.8900 5.7950 0.8900
                 5.7950 1.3300 6.2750 1.3300 6.2750 1.1900 6.3950 1.1900 ;
        POLYGON  6.0350 1.2100 5.9150 1.2100 5.9150 0.5300 4.4450 0.5300 4.4450 1.1600 3.7150 1.1600
                 3.7150 1.7250 3.3400 1.7250 3.3400 2.0100 2.9150 2.0100 2.9150 1.8900 3.2200 1.8900
                 3.2200 1.6050 3.5950 1.6050 3.5950 0.9000 3.2550 0.9000 3.2550 0.8600 3.1350 0.8600
                 3.1350 0.7400 3.3750 0.7400 3.3750 0.7800 3.7150 0.7800 3.7150 1.0400 4.3250 1.0400
                 4.3250 0.4100 6.0350 0.4100 ;
        POLYGON  4.3750 1.9650 3.5800 1.9650 3.5800 2.2500 2.6650 2.2500 2.6650 1.9700 2.4150 1.9700
                 2.4150 1.9650 1.7400 1.9650 1.7400 1.9700 1.4750 1.9700 1.4750 2.0900 1.3550 2.0900
                 1.3550 1.9700 1.2750 1.9700 1.2750 0.6600 1.3950 0.6600 1.3950 1.8500 1.6200 1.8500
                 1.6200 1.8450 2.5350 1.8450 2.5350 1.8500 2.7850 1.8500 2.7850 2.1300 3.4600 2.1300
                 3.4600 1.8450 4.2550 1.8450 4.2550 1.3300 4.3750 1.3300 ;
        POLYGON  3.4750 1.2600 3.3550 1.2600 3.3550 1.1700 2.9350 1.1700 2.9350 1.7300 2.8150 1.7300
                 2.8150 1.1700 1.9950 1.1700 1.9950 1.1800 1.7550 1.1800 1.7550 1.0500 3.3550 1.0500
                 3.3550 1.0200 3.4750 1.0200 ;
        POLYGON  3.0350 0.6200 1.6350 0.6200 1.6350 1.7250 1.5150 1.7250 1.5150 0.5400 0.9750 0.5400
                 0.9750 1.0800 0.2400 1.0800 0.2400 1.8500 0.3550 1.8500 0.3550 2.0900 0.2350 2.0900
                 0.2350 1.9700 0.1200 1.9700 0.1200 0.7800 0.1350 0.7800 0.1350 0.6600 0.2550 0.6600
                 0.2550 0.9600 0.8550 0.9600 0.8550 0.4200 0.9950 0.4200 0.9950 0.4000 1.2350 0.4000
                 1.2350 0.4200 1.6350 0.4200 1.6350 0.5000 2.9150 0.5000 2.9150 0.3600 3.0350 0.3600 ;
    END
END MXI4X4

MACRO MXI4X2
    CLASS CORE ;
    FOREIGN MXI4X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4200 1.1450 4.5700 1.4350 ;
        RECT  4.3100 1.1400 4.4300 1.4200 ;
        END
    END D
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5550 1.2300 7.8150 1.3800 ;
        RECT  7.5550 1.1400 7.7950 1.3800 ;
        RECT  7.4750 1.3800 7.6300 1.5000 ;
        RECT  7.2100 1.5550 7.5950 1.6750 ;
        RECT  7.4750 1.3800 7.5950 1.6750 ;
        RECT  7.5100 1.2600 7.5950 1.6750 ;
        RECT  4.9300 1.9600 7.3300 2.0800 ;
        RECT  7.2100 1.5550 7.3300 2.0800 ;
        RECT  5.0100 1.2400 5.1300 1.4800 ;
        RECT  4.9300 1.3600 5.0500 2.0800 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.5000 1.0300 1.6300 ;
        RECT  0.6500 1.4650 0.8000 1.7500 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.5400 2.4250 1.7800 ;
        RECT  2.0450 1.5200 2.3050 1.7800 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3288  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.8267  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 1.1600 1.3300 1.4000 ;
        RECT  0.3600 1.2250 1.3300 1.3450 ;
        RECT  0.4100 1.2250 0.5300 1.4650 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.5400 2.9300 1.7700 ;
        RECT  2.6250 1.5200 2.8850 1.7700 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9700 1.1750 7.1800 1.4350 ;
        RECT  6.9700 0.7400 7.0900 1.8400 ;
        RECT  6.8500 0.7400 7.0900 0.8600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.4500 -0.1800 7.5700 0.7800 ;
        RECT  6.1300 0.6000 6.3700 0.7200 ;
        RECT  6.1300 -0.1800 6.2500 0.7200 ;
        RECT  4.3300 -0.1800 4.4500 0.7800 ;
        RECT  2.4900 -0.1800 2.6100 0.6800 ;
        RECT  0.6500 -0.1800 0.7700 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.4500 2.0600 7.5700 2.7900 ;
        RECT  6.4900 2.2000 6.6100 2.7900 ;
        RECT  4.3900 2.2800 4.6300 2.7900 ;
        RECT  2.4900 2.1400 2.6100 2.7900 ;
        RECT  0.5900 1.9600 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.0550 1.6200 7.7500 1.6200 7.7500 1.5000 7.9350 1.5000 7.9350 1.0200 7.2100 1.0200
                 7.2100 0.6200 6.6100 0.6200 6.6100 1.6000 5.4100 1.6000 5.4100 1.1200 4.9300 1.1200
                 4.9300 1.0600 4.8100 1.0600 4.8100 0.9400 5.0500 0.9400 5.0500 1.0000 5.5300 1.0000
                 5.5300 1.4800 6.4900 1.4800 6.4900 0.5000 7.3300 0.5000 7.3300 0.9000 7.9300 0.9000
                 7.9300 0.6600 8.0500 0.6600 8.0500 0.7800 8.0550 0.7800 ;
        POLYGON  6.8500 1.8400 5.1700 1.8400 5.1700 1.6000 5.2900 1.6000 5.2900 1.7200 6.7300 1.7200
                 6.7300 1.1800 6.8500 1.1800 ;
        POLYGON  6.3700 1.3600 5.6500 1.3600 5.6500 0.8800 5.1700 0.8800 5.1700 0.7200 4.9700 0.7200
                 4.9700 0.6000 5.2900 0.6000 5.2900 0.7600 5.7700 0.7600 5.7700 1.2400 6.3700 1.2400 ;
        POLYGON  6.1300 1.0400 5.8900 1.0400 5.8900 0.4800 4.6900 0.4800 4.6900 1.0200 4.1900 1.0200
                 4.1900 1.9200 3.8100 1.9200 3.8100 2.0000 3.5700 2.0000 3.5700 1.8800 3.6900 1.8800
                 3.6900 1.8000 4.0700 1.8000 4.0700 0.8800 3.6300 0.8800 3.6300 0.6200 3.7500 0.6200
                 3.7500 0.7600 4.1900 0.7600 4.1900 0.9000 4.5700 0.9000 4.5700 0.3600 6.0100 0.3600
                 6.0100 0.9200 6.1300 0.9200 ;
        POLYGON  4.8100 2.1600 4.0500 2.1600 4.0500 2.2400 3.3050 2.2400 3.3050 2.0200 1.5700 2.0200
                 1.5700 2.0800 1.4500 2.0800 1.4500 0.6200 1.5700 0.6200 1.5700 1.9000 3.4250 1.9000
                 3.4250 2.1200 3.9300 2.1200 3.9300 2.0400 4.6900 2.0400 4.6900 1.2400 4.8100 1.2400 ;
        POLYGON  3.9500 1.1200 3.8300 1.1200 3.8300 1.4000 3.1900 1.4000 3.1900 1.7200 3.0700 1.7200
                 3.0700 1.4000 1.9300 1.4000 1.9300 1.1600 2.0500 1.1600 2.0500 1.2800 3.7100 1.2800
                 3.7100 1.0000 3.9500 1.0000 ;
        POLYGON  3.9500 1.6800 3.7100 1.6800 3.7100 1.6400 3.3500 1.6400 3.3500 1.5200 3.8300 1.5200
                 3.8300 1.5600 3.9500 1.5600 ;
        RECT  2.9900 1.0400 3.5900 1.1600 ;
        POLYGON  3.2300 0.4800 3.1100 0.4800 3.1100 0.9200 2.1950 0.9200 2.1950 0.5000 1.8100 0.5000
                 1.8100 1.7600 1.6900 1.7600 1.6900 0.5000 1.0150 0.5000 1.0150 1.0400 0.2400 1.0400
                 0.2400 1.5550 0.2900 1.5550 0.2900 2.0800 0.1700 2.0800 0.1700 1.6750 0.1200 1.6750
                 0.1200 0.8000 0.1700 0.8000 0.1700 0.6800 0.2900 0.6800 0.2900 0.9200 0.8950 0.9200
                 0.8950 0.3800 1.1600 0.3800 1.1600 0.3600 1.4000 0.3600 1.4000 0.3800 2.3150 0.3800
                 2.3150 0.8000 2.9900 0.8000 2.9900 0.3600 3.2300 0.3600 ;
    END
END MXI4X2

MACRO MXI4X1
    CLASS CORE ;
    FOREIGN MXI4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4650 0.4400 2.5850 1.0400 ;
        RECT  2.4450 0.9200 2.5650 1.5300 ;
        RECT  1.8200 0.4400 2.5850 0.5600 ;
        RECT  1.9650 0.3600 2.2050 0.5600 ;
        RECT  0.7750 0.4800 1.9400 0.6000 ;
        RECT  0.7750 0.4800 0.8950 1.2400 ;
        RECT  0.6500 0.5950 0.8950 0.8550 ;
        END
    END S1
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9750 1.2650 3.4250 1.3900 ;
        RECT  2.9150 1.2300 3.3450 1.3850 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0750 1.5200 4.5250 1.6700 ;
        RECT  4.4050 1.4300 4.5250 1.6700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6450 1.4800 4.9600 1.7050 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8150 1.5250 6.2050 1.7050 ;
        RECT  5.8150 1.5000 6.0750 1.7050 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.1560  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        ANTENNAMAXAREACAR 0.8667  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7450 1.2400 6.5450 1.3600 ;
        RECT  6.1050 1.2300 6.3650 1.3800 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6600 0.2550 2.0600 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  6.2250 -0.1800 6.3450 0.3800 ;
        RECT  4.8250 -0.1800 4.9450 0.8300 ;
        RECT  3.1050 -0.1800 3.2250 0.8600 ;
        RECT  1.4050 -0.1800 1.6450 0.3600 ;
        RECT  0.5550 -0.1800 0.7950 0.3200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  6.1450 1.9400 6.2650 2.7900 ;
        RECT  4.5400 2.0650 4.6600 2.7900 ;
        RECT  4.4200 2.0650 4.6600 2.1850 ;
        RECT  2.9850 2.2200 3.2250 2.7900 ;
        RECT  1.2250 1.9100 1.4650 2.0300 ;
        RECT  1.2250 1.9100 1.3450 2.7900 ;
        RECT  0.4950 1.8800 0.7350 2.0000 ;
        RECT  0.4950 1.8800 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.8250 0.9000 6.7850 0.9000 6.7850 1.6000 6.6850 1.6000 6.6850 2.0600 6.5650 2.0600
                 6.5650 1.4800 6.6650 1.4800 6.6650 0.7800 6.7050 0.7800 6.7050 0.6200 5.9100 0.6200
                 5.9100 0.5800 5.3450 0.5800 5.3450 0.9500 5.3850 0.9500 5.3850 1.7400 5.2650 1.7400
                 5.2650 1.0700 4.3900 1.0700 4.3900 0.5600 3.7050 0.5600 3.7050 1.6200 3.5850 1.6200
                 3.5850 0.4400 4.0050 0.4400 4.0050 0.3600 4.2450 0.3600 4.2450 0.4400 4.5100 0.4400
                 4.5100 0.9500 5.2250 0.9500 5.2250 0.4600 5.6250 0.4600 5.6250 0.3600 5.8650 0.3600
                 5.8650 0.4600 6.0300 0.4600 6.0300 0.5000 6.8250 0.5000 ;
        POLYGON  5.7050 0.8200 5.6250 0.8200 5.6250 2.0600 5.5050 2.0600 5.5050 1.9800 4.9750 1.9800
                 4.9750 1.9450 4.3000 1.9450 4.3000 2.2500 3.3850 2.2500 3.3850 2.1000 2.8650 2.1000
                 2.8650 2.2500 2.6250 2.2500 2.6250 2.1300 2.7450 2.1300 2.7450 1.9800 3.5050 1.9800
                 3.5050 2.1300 4.1800 2.1300 4.1800 1.8250 5.0950 1.8250 5.0950 1.8600 5.5050 1.8600
                 5.5050 0.8200 5.4650 0.8200 5.4650 0.7000 5.7050 0.7000 ;
        POLYGON  5.1450 1.3600 4.9050 1.3600 4.9050 1.3100 4.1850 1.3100 4.1850 1.3800 4.0650 1.3800
                 4.0650 1.1400 4.1850 1.1400 4.1850 1.1900 5.1450 1.1900 ;
        POLYGON  4.1050 0.8000 3.9450 0.8000 3.9450 1.8900 3.8650 1.8900 3.8650 2.0100 3.7450 2.0100
                 3.7450 1.8600 2.6250 1.8600 2.6250 1.9900 2.5050 1.9900 2.5050 2.1100 1.8250 2.1100
                 1.8250 2.2500 1.5850 2.2500 1.5850 2.1300 1.7050 2.1300 1.7050 1.9900 2.3850 1.9900
                 2.3850 1.8700 2.5050 1.8700 2.5050 1.7400 3.8250 1.7400 3.8250 0.6800 4.1050 0.6800 ;
        POLYGON  2.3450 0.8000 2.3250 0.8000 2.3250 1.7500 2.2650 1.7500 2.2650 1.8700 2.1450 1.8700
                 2.1450 1.7600 0.4150 1.7600 0.4150 1.0200 0.5350 1.0200 0.5350 1.6400 2.1450 1.6400
                 2.1450 1.6300 2.2050 1.6300 2.2050 0.8000 2.1050 0.8000 2.1050 0.6800 2.3450 0.6800 ;
        POLYGON  2.0850 1.5100 1.2150 1.5100 1.2150 1.5200 0.9750 1.5200 0.9750 1.4000 1.0950 1.4000
                 1.0950 0.8400 1.0150 0.8400 1.0150 0.7200 1.2550 0.7200 1.2550 0.8400 1.2150 0.8400
                 1.2150 1.3900 1.9650 1.3900 1.9650 1.2700 2.0850 1.2700 ;
    END
END MXI4X1

MACRO MXI3XL
    CLASS CORE ;
    FOREIGN MXI3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3350 1.4650 1.5750 1.5850 ;
        RECT  0.3050 1.5200 1.4550 1.6200 ;
        RECT  0.3550 1.5000 1.5750 1.5850 ;
        RECT  0.3050 1.5200 0.5650 1.6700 ;
        RECT  0.3550 1.3800 0.4750 1.6700 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2300 1.1150 1.3500 ;
        RECT  0.5950 1.2300 0.8550 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3150 1.3950 2.5400 1.7250 ;
        END
    END B
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5150 1.4200 4.4750 1.5400 ;
        RECT  3.5150 1.2300 3.7550 1.5400 ;
        RECT  3.5150 1.1800 3.6350 1.5400 ;
        RECT  3.4950 1.2300 3.7550 1.3800 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9650 1.1750 5.1750 1.4350 ;
        RECT  4.9650 1.0400 5.1500 1.4350 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6650 0.6800 5.7850 1.6000 ;
        RECT  5.5800 0.8850 5.7850 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.2450 -0.1800 5.3650 0.9200 ;
        RECT  3.9550 0.7000 4.1950 0.8200 ;
        RECT  3.9550 -0.1800 4.0750 0.8200 ;
        RECT  2.2550 0.7000 2.4950 0.8200 ;
        RECT  2.2550 -0.1800 2.3750 0.8200 ;
        RECT  0.7550 -0.1800 0.8750 0.8700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1250 2.1000 5.3650 2.2200 ;
        RECT  5.1250 2.1000 5.2450 2.7900 ;
        RECT  3.6950 2.2650 3.9350 2.7900 ;
        RECT  2.3150 1.8450 2.4350 2.7900 ;
        RECT  0.8750 1.8450 0.9950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7050 1.9800 5.0050 1.9800 5.0050 2.1450 3.8300 2.1450 3.8300 2.1000 3.0350 2.1000
                 3.0350 1.8600 2.8550 1.8600 2.8550 0.7000 3.1350 0.7000 3.1350 0.8200 2.9750 0.8200
                 2.9750 1.7400 3.1550 1.7400 3.1550 1.9800 3.9500 1.9800 3.9500 2.0250 4.8850 2.0250
                 4.8850 1.8600 5.7050 1.8600 ;
        POLYGON  4.9450 0.9200 4.8450 0.9200 4.8450 1.3000 4.8250 1.3000 4.8250 1.6000 4.7050 1.6000
                 4.7050 1.3000 3.8750 1.3000 3.8750 1.1800 4.7250 1.1800 4.7250 0.8000 4.8250 0.8000
                 4.8250 0.6800 4.9450 0.6800 ;
        POLYGON  4.5550 1.0600 3.3750 1.0600 3.3750 1.5000 3.3950 1.5000 3.3950 1.6650 4.2950 1.6650
                 4.2950 1.7850 4.4150 1.7850 4.4150 1.9050 4.1750 1.9050 4.1750 1.7850 3.2750 1.7850
                 3.2750 1.6200 3.2150 1.6200 3.2150 1.5850 3.0950 1.5850 3.0950 1.4650 3.2550 1.4650
                 3.2550 0.5800 2.8550 0.5800 2.8550 0.4800 2.7350 0.4800 2.7350 0.3600 2.9750 0.3600
                 2.9750 0.4600 3.5050 0.4600 3.5050 0.9400 4.4350 0.9400 4.4350 0.6400 4.5550 0.6400 ;
        POLYGON  2.5950 1.2750 2.4750 1.2750 2.4750 1.2650 2.1950 1.2650 2.1950 1.8650 1.8550 1.8650
                 1.8550 1.9050 1.6150 1.9050 1.6150 1.7850 1.7350 1.7850 1.7350 1.7450 2.0750 1.7450
                 2.0750 1.2650 2.0150 1.2650 2.0150 0.8200 1.3950 0.8200 1.3950 0.7000 2.1350 0.7000
                 2.1350 1.1450 2.4750 1.1450 2.4750 1.0350 2.5950 1.0350 ;
        POLYGON  1.9550 1.6250 1.8350 1.6250 1.8350 1.5050 1.6950 1.5050 1.6950 1.1600 1.2350 1.1600
                 1.2350 1.1100 0.1850 1.1100 0.1850 1.7900 0.5750 1.7900 0.5750 2.0300 0.4550 2.0300
                 0.4550 1.9100 0.0650 1.9100 0.0650 0.8700 0.2750 0.8700 0.2750 0.6400 0.3950 0.6400
                 0.3950 0.9900 1.8150 0.9900 1.8150 1.3850 1.9550 1.3850 ;
    END
END MXI3XL

MACRO MXI3X4
    CLASS CORE ;
    FOREIGN MXI3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2550 1.0000 0.3750 1.2400 ;
        RECT  0.0700 1.0000 0.3750 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2850 1.4100 2.5650 1.5300 ;
        RECT  2.2850 1.0900 2.4050 1.5300 ;
        RECT  1.7250 1.0900 2.4050 1.2100 ;
        RECT  1.8050 0.8850 1.9600 1.2100 ;
        RECT  1.7250 1.0900 1.8450 1.3400 ;
        RECT  1.2450 1.1800 1.9250 1.3000 ;
        RECT  1.1250 1.3000 1.3650 1.4200 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6850 1.2000 4.8050 1.4400 ;
        RECT  4.4200 1.2000 4.8050 1.4350 ;
        RECT  4.4200 1.1750 4.5700 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9650 1.2300 6.3650 1.4800 ;
        RECT  6.1050 1.2100 6.3650 1.4800 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3450 0.9700 6.5250 1.0900 ;
        RECT  5.7250 0.9400 6.0750 1.0900 ;
        RECT  5.7250 0.9300 5.8450 1.1700 ;
        RECT  5.1650 1.3800 5.4650 1.5000 ;
        RECT  5.3450 0.9700 5.4650 1.5000 ;
        RECT  5.1650 1.3800 5.2850 1.6200 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4450 0.6900 4.6450 0.8100 ;
        RECT  4.1850 1.5550 4.3050 2.2100 ;
        RECT  4.1800 0.6900 4.3000 1.6750 ;
        RECT  3.5250 1.3200 4.3000 1.4400 ;
        RECT  3.5500 1.1750 3.7000 1.4400 ;
        RECT  3.3450 1.4600 3.6450 1.5800 ;
        RECT  3.5250 1.3200 3.6450 1.5800 ;
        RECT  3.3450 1.4600 3.4650 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  6.2850 -0.1800 6.4050 0.8100 ;
        RECT  4.8850 -0.1800 5.1250 0.3300 ;
        RECT  3.9250 -0.1800 4.1650 0.3300 ;
        RECT  2.9650 -0.1800 3.0850 0.6800 ;
        RECT  1.4650 -0.1800 1.5850 0.6800 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  6.0850 1.8400 6.2050 2.7900 ;
        RECT  4.6050 1.5600 4.7250 2.7900 ;
        RECT  3.7650 1.5600 3.8850 2.7900 ;
        RECT  2.9250 1.5600 3.0450 2.7900 ;
        RECT  1.5650 1.7800 1.6850 2.7900 ;
        RECT  0.1350 1.4600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.8250 0.8100 6.7650 0.8100 6.7650 1.8400 6.6250 1.8400 6.6250 1.9600 6.5050 1.9600
                 6.5050 1.7200 5.5850 1.7200 5.5850 1.4000 5.7050 1.4000 5.7050 1.6000 6.6450 1.6000
                 6.6450 0.6900 6.7050 0.6900 6.7050 0.5700 6.8250 0.5700 ;
        POLYGON  5.7650 0.8100 5.6450 0.8100 5.6450 0.6900 5.0450 0.6900 5.0450 1.7400 5.4450 1.7400
                 5.4450 1.9800 5.3250 1.9800 5.3250 1.8600 4.9250 1.8600 4.9250 0.6900 4.7950 0.6900
                 4.7950 0.5700 3.3250 0.5700 3.3250 0.9200 3.0050 0.9200 3.0050 1.0400 2.7650 1.0400
                 2.7650 0.9200 2.8850 0.9200 2.8850 0.8000 3.2050 0.8000 3.2050 0.4500 4.9150 0.4500
                 4.9150 0.5700 5.7650 0.5700 ;
        POLYGON  3.4050 1.3400 2.8050 1.3400 2.8050 1.7700 2.4050 1.7700 2.4050 1.8100 2.3450 1.8100
                 2.3450 2.2100 2.2250 2.2100 2.2250 1.6900 2.2850 1.6900 2.2850 1.6500 2.6850 1.6500
                 2.6850 1.2800 2.5250 1.2800 2.5250 0.7800 2.1050 0.7800 2.1050 0.5400 2.2250 0.5400
                 2.2250 0.6600 2.6450 0.6600 2.6450 1.1600 2.8050 1.1600 2.8050 1.2200 3.4050 1.2200 ;
        POLYGON  2.1650 1.5700 2.1050 1.5700 2.1050 1.6600 1.1450 1.6600 1.1450 1.9300 1.0250 1.9300
                 1.0250 1.7800 0.8850 1.7800 0.8850 0.7200 0.8650 0.7200 0.8650 0.6000 1.1050 0.6000
                 1.1050 0.7200 1.0050 0.7200 1.0050 1.5400 1.9850 1.5400 1.9850 1.4500 2.0450 1.4500
                 2.0450 1.3300 2.1650 1.3300 ;
        POLYGON  1.5850 1.0600 1.3450 1.0600 1.3450 0.9200 1.2250 0.9200 1.2250 0.4800 0.6550 0.4800
                 0.6550 0.8000 0.6750 0.8000 0.6750 1.5800 0.5550 1.5800 0.5550 0.9200 0.5350 0.9200
                 0.5350 0.3600 1.3450 0.3600 1.3450 0.8000 1.4650 0.8000 1.4650 0.9400 1.5850 0.9400 ;
    END
END MXI3X4

MACRO MXI3X2
    CLASS CORE ;
    FOREIGN MXI3X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.3950 1.2950 ;
        RECT  0.2750 1.0550 0.3950 1.2950 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.5200 2.9500 1.6400 ;
        RECT  2.8300 1.2400 2.9500 1.6400 ;
        RECT  2.2900 1.0200 2.4100 1.6400 ;
        RECT  2.0450 1.5200 2.3050 1.6700 ;
        RECT  1.2300 1.2600 1.3500 1.6400 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1300 1.1750 4.5300 1.2950 ;
        RECT  4.4100 1.0550 4.5300 1.2950 ;
        RECT  4.1300 1.1750 4.2800 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8700 1.1100 6.0500 1.5000 ;
        RECT  5.9300 1.1000 6.0500 1.5000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3950 0.9400 6.6550 1.0900 ;
        RECT  5.1100 0.8600 6.5150 0.9800 ;
        RECT  6.2900 0.9400 6.6550 1.0600 ;
        RECT  5.6100 0.8400 5.7300 1.0800 ;
        RECT  4.8900 1.4000 5.2300 1.5200 ;
        RECT  5.1100 0.8600 5.2300 1.5200 ;
        RECT  4.8900 1.4000 5.0100 1.6400 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8100 0.7400 4.0500 0.8600 ;
        RECT  3.8700 0.7400 3.9900 2.2100 ;
        RECT  3.8400 1.1750 3.9900 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  6.0900 -0.1800 6.2100 0.7400 ;
        RECT  4.2900 -0.1800 4.5300 0.3800 ;
        RECT  3.3300 -0.1800 3.5700 0.3800 ;
        RECT  1.4300 -0.1800 1.5500 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  5.9900 1.8600 6.1100 2.7900 ;
        RECT  4.2900 1.5600 4.4100 2.7900 ;
        RECT  3.4500 1.5800 3.5700 2.7900 ;
        RECT  1.4300 2.2200 1.5500 2.7900 ;
        RECT  0.1350 1.5550 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.8950 1.8600 6.5300 1.8600 6.5300 1.9800 6.4100 1.9800 6.4100 1.7400 5.3500 1.7400
                 5.3500 1.4200 5.4700 1.4200 5.4700 1.6200 6.7750 1.6200 6.7750 0.7400 6.5100 0.7400
                 6.5100 0.5000 6.6300 0.5000 6.6300 0.6200 6.8950 0.6200 ;
        POLYGON  5.4900 0.7400 5.3700 0.7400 5.3700 0.6200 4.7700 0.6200 4.7700 1.7600 5.1100 1.7600
                 5.1100 1.8000 5.2300 1.8000 5.2300 1.9200 4.9900 1.9200 4.9900 1.8800 4.6500 1.8800
                 4.6500 0.6200 3.0900 0.6200 3.0900 0.5400 2.9700 0.5400 2.9700 0.4200 3.2100 0.4200
                 3.2100 0.5000 5.4900 0.5000 ;
        POLYGON  3.7100 1.2400 3.5900 1.2400 3.5900 1.1200 3.1900 1.1200 3.1900 1.8800 2.6100 1.8800
                 2.6100 1.7600 3.0700 1.7600 3.0700 1.1200 2.5300 1.1200 2.5300 0.6800 2.6500 0.6800
                 2.6500 1.0000 3.7100 1.0000 ;
        POLYGON  2.0900 1.4000 1.9700 1.4000 1.9700 1.1400 1.0700 1.1400 1.0700 1.8200 0.9500 1.8200
                 0.9500 0.6800 1.0700 0.6800 1.0700 1.0200 2.0900 1.0200 ;
        POLYGON  1.9500 0.5400 1.8300 0.5400 1.8300 0.6200 1.1900 0.6200 1.1900 0.5600 0.7800 0.5600
                 0.7800 0.6800 0.6750 0.6800 0.6750 1.6750 0.5550 1.6750 0.5550 0.5600 0.6600 0.5600
                 0.6600 0.4400 1.3100 0.4400 1.3100 0.5000 1.7100 0.5000 1.7100 0.4200 1.9500 0.4200 ;
    END
END MXI3X2

MACRO MXI3X1
    CLASS CORE ;
    FOREIGN MXI3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.5200 1.4550 1.6400 ;
        RECT  1.3350 1.3600 1.4550 1.6400 ;
        RECT  0.3050 1.5200 0.5650 1.6700 ;
        RECT  0.3550 1.3400 0.4750 1.6700 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2100 1.0350 1.3650 ;
        RECT  0.5950 1.2100 0.8550 1.4000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3350 1.5000 2.5950 1.6700 ;
        RECT  2.2550 1.3400 2.3750 1.6200 ;
        END
    END B
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4550 1.4000 4.4750 1.5200 ;
        RECT  3.4550 1.2300 3.7550 1.5200 ;
        RECT  3.4550 1.1600 3.6950 1.5200 ;
        END
    END S1
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 0.9000 5.2050 1.1150 ;
        RECT  4.9650 0.9000 5.0850 1.2800 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6650 0.6800 5.7850 1.9900 ;
        RECT  5.5800 0.8850 5.7850 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.2450 -0.1800 5.3650 0.7800 ;
        RECT  3.9550 0.6800 4.1950 0.8000 ;
        RECT  3.9550 -0.1800 4.0750 0.8000 ;
        RECT  2.2750 -0.1800 2.3950 0.8600 ;
        RECT  0.6550 0.6800 0.8950 0.8000 ;
        RECT  0.6550 -0.1800 0.7750 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1250 1.8800 5.3650 2.0000 ;
        RECT  5.1250 1.8800 5.2450 2.7900 ;
        RECT  3.6950 2.2200 3.9350 2.7900 ;
        RECT  2.3350 1.8000 2.4550 2.7900 ;
        RECT  0.7950 1.8000 0.9150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.4600 1.5200 5.2150 1.5200 5.2150 1.7600 4.9500 1.7600 4.9500 2.1000 2.9750 2.1000
                 2.9750 1.8600 2.8550 1.8600 2.8550 0.6800 3.0950 0.6800 3.0950 0.8000 2.9750 0.8000
                 2.9750 1.7400 3.0950 1.7400 3.0950 1.9800 4.8300 1.9800 4.8300 1.6400 5.0950 1.6400
                 5.0950 1.4000 5.3400 1.4000 5.3400 1.0200 5.4600 1.0200 ;
        POLYGON  4.9450 0.7800 4.7950 0.7800 4.7950 1.2800 4.7650 1.2800 4.7650 1.4000 4.8850 1.4000
                 4.8850 1.5200 4.6450 1.5200 4.6450 1.2800 3.8750 1.2800 3.8750 1.1600 4.6750 1.1600
                 4.6750 0.6600 4.8250 0.6600 4.8250 0.5400 4.9450 0.5400 ;
        POLYGON  4.5550 1.0400 3.6400 1.0400 3.6400 0.5600 3.3350 0.5600 3.3350 1.6400 4.2950 1.6400
                 4.2950 1.7400 4.4150 1.7400 4.4150 1.8600 4.1750 1.8600 4.1750 1.7600 3.2150 1.7600
                 3.2150 1.5400 3.0950 1.5400 3.0950 1.4200 3.2150 1.4200 3.2150 0.5600 3.1000 0.5600
                 3.1000 0.4800 2.7150 0.4800 2.7150 0.3600 3.2200 0.3600 3.2200 0.4400 3.7600 0.4400
                 3.7600 0.9200 4.4350 0.9200 4.4350 0.6200 4.5550 0.6200 ;
        POLYGON  2.5550 1.2200 2.1350 1.2200 2.1350 1.8200 1.7950 1.8200 1.7950 1.8800 1.5550 1.8800
                 1.5550 1.7600 1.6750 1.7600 1.6750 1.7000 2.0150 1.7000 2.0150 1.2200 1.8150 1.2200
                 1.8150 0.8000 1.2950 0.8000 1.2950 0.6800 1.9350 0.6800 1.9350 1.1000 2.4350 1.1000
                 2.4350 0.9800 2.5550 0.9800 ;
        POLYGON  1.8950 1.5800 1.7750 1.5800 1.7750 1.4600 1.5750 1.4600 1.5750 1.1200 1.1550 1.1200
                 1.1550 1.0900 0.1850 1.0900 0.1850 1.7900 0.4950 1.7900 0.4950 2.0300 0.3750 2.0300
                 0.3750 1.9100 0.0650 1.9100 0.0650 0.7400 0.2950 0.7400 0.2950 0.6200 0.4150 0.6200
                 0.4150 0.9700 1.6950 0.9700 1.6950 1.3400 1.8950 1.3400 ;
    END
END MXI3X1

MACRO MXI2XL
    CLASS CORE ;
    FOREIGN MXI2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1500 1.2650 0.2700 1.5950 ;
        RECT  0.0700 1.1000 0.2200 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2200 1.4400 1.4000 1.8500 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.2000 1.7400 1.4400 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.5500 1.2000 1.6700 1.7250 ;
        RECT  0.8700 1.2000 1.7400 1.3200 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1920  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.7200 0.9600 0.8400 ;
        RECT  0.7800 1.8900 0.9000 2.1300 ;
        RECT  0.3900 1.8900 0.9000 2.0100 ;
        RECT  0.3900 0.7200 0.5100 2.0100 ;
        RECT  0.3600 0.8850 0.5100 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3700 0.7200 1.6100 0.8400 ;
        RECT  1.3700 -0.1800 1.4900 0.8400 ;
        RECT  0.1350 -0.1800 0.2550 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.4200 1.9700 1.5400 2.7900 ;
        RECT  0.1400 1.9700 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9800 1.6800 1.9600 1.6800 1.9600 2.0900 1.8400 2.0900 1.8400 1.5600 1.8600 1.5600
                 1.8600 1.0800 0.7500 1.0800 0.7500 1.4400 1.0400 1.4400 1.0400 1.7700 0.9200 1.7700
                 0.9200 1.5600 0.6300 1.5600 0.6300 0.9600 1.0800 0.9600 1.0800 0.6000 0.6800 0.6000
                 0.6800 0.5000 0.5600 0.5000 0.5600 0.3800 0.8000 0.3800 0.8000 0.4800 1.2500 0.4800
                 1.2500 0.9600 1.8500 0.9600 1.8500 0.6600 1.9700 0.6600 1.9700 0.7800 1.9800 0.7800 ;
    END
END MXI2XL

MACRO MXI2X8
    CLASS CORE ;
    FOREIGN MXI2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.5550 1.2700 1.6750 ;
        RECT  1.1500 1.4050 1.2700 1.6750 ;
        RECT  0.4100 1.5050 0.5300 1.7450 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.9500 1.4150 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.9500 1.1750 2.2500 1.4050 ;
        RECT  1.9500 1.1650 2.0700 1.4050 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7900 1.2200 5.9100 2.2000 ;
        RECT  4.1700 0.7900 5.9100 0.9100 ;
        RECT  5.7900 0.6700 5.9100 0.9100 ;
        RECT  3.2600 1.2200 5.9100 1.3400 ;
        RECT  5.4800 0.7900 5.6000 1.3400 ;
        RECT  4.8900 0.7400 5.1300 0.9100 ;
        RECT  4.9500 1.2200 5.0700 2.2000 ;
        RECT  4.0500 0.7400 4.2900 0.8600 ;
        RECT  4.1100 1.2200 4.2300 2.2050 ;
        RECT  3.2600 1.1750 3.4100 1.4350 ;
        RECT  3.2700 0.6800 3.3900 2.2050 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.3700 -0.1800 5.4900 0.6700 ;
        RECT  4.5300 -0.1800 4.6500 0.6700 ;
        RECT  3.6900 -0.1800 3.8100 0.6700 ;
        RECT  2.8500 -0.1800 2.9700 0.7300 ;
        RECT  2.0100 -0.1800 2.1300 0.8050 ;
        RECT  0.6700 -0.1800 0.7900 0.8050 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.3700 1.4600 5.4900 2.7900 ;
        RECT  4.5300 1.4600 4.6500 2.7900 ;
        RECT  3.6900 1.4600 3.8100 2.7900 ;
        RECT  2.8500 1.5550 2.9700 2.7900 ;
        RECT  2.0100 1.5550 2.1300 2.7900 ;
        RECT  0.6700 1.9650 0.7900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1400 1.3200 2.7300 1.3200 2.7300 1.6750 2.5500 1.6750 2.5500 2.2050 2.4300 2.2050
                 2.4300 1.5550 2.6100 1.5550 2.6100 0.8050 2.4300 0.8050 2.4300 0.5650 2.5500 0.5650
                 2.5500 0.6850 2.7300 0.6850 2.7300 1.2000 3.1400 1.2000 ;
        POLYGON  2.4900 1.2400 2.3700 1.2400 2.3700 1.0450 1.8300 1.0450 1.8300 1.9850 1.4900 1.9850
                 1.4900 2.0250 1.2500 2.0250 1.2500 1.9050 1.3700 1.9050 1.3700 1.8650 1.7100 1.8650
                 1.7100 1.0450 1.3900 1.0450 1.3900 0.8050 1.3100 0.8050 1.3100 0.5650 1.4300 0.5650
                 1.4300 0.6850 1.5100 0.6850 1.5100 0.9250 2.4900 0.9250 ;
        POLYGON  1.5900 1.7450 1.4700 1.7450 1.4700 1.2850 1.1500 1.2850 1.1500 1.0550 0.2400 1.0550
                 0.2400 1.8450 0.2900 1.8450 0.2900 2.0850 0.1700 2.0850 0.1700 1.9650 0.1200 1.9650
                 0.1200 0.6850 0.2500 0.6850 0.2500 0.5650 0.3700 0.5650 0.3700 0.8050 0.2400 0.8050
                 0.2400 0.9350 1.1500 0.9350 1.1500 0.9250 1.2700 0.9250 1.2700 1.1650 1.5900 1.1650 ;
    END
END MXI2X8

MACRO MXI2X6
    CLASS CORE ;
    FOREIGN MXI2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4100 1.5550 1.1900 1.6750 ;
        RECT  1.0700 1.0950 1.1900 1.6750 ;
        RECT  0.4100 1.3150 0.5300 1.6750 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0950 0.8700 1.4200 ;
        RECT  0.6500 1.1050 0.8350 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.8900 1.1750 2.2500 1.4150 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0300 0.4050 5.1500 1.0400 ;
        RECT  4.9500 1.1900 5.0700 2.2100 ;
        RECT  4.8500 0.9200 5.1500 1.0400 ;
        RECT  4.1900 1.0400 4.9700 1.3100 ;
        RECT  4.1900 0.4050 4.3100 1.3100 ;
        RECT  4.1100 1.1900 4.2300 2.2100 ;
        RECT  3.5500 1.1900 5.0700 1.3100 ;
        RECT  3.5500 1.1750 3.7000 1.4350 ;
        RECT  3.2900 1.0700 3.6700 1.1900 ;
        RECT  3.2700 1.3100 3.7000 1.4300 ;
        RECT  3.2900 0.4000 3.4100 1.1900 ;
        RECT  3.2700 1.3100 3.3900 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.6100 -0.1800 4.7300 0.9200 ;
        RECT  3.7700 -0.1800 3.8900 0.9200 ;
        RECT  2.8700 -0.1800 2.9900 0.8450 ;
        RECT  2.0300 -0.1800 2.1500 0.6550 ;
        RECT  0.7500 -0.1800 0.8700 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.5300 1.4300 4.6500 2.7900 ;
        RECT  3.6900 1.5550 3.8100 2.7900 ;
        RECT  2.8500 1.5600 2.9700 2.7900 ;
        RECT  2.0100 1.6750 2.1300 2.7900 ;
        RECT  0.6700 1.7950 0.7900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1500 1.2600 2.7300 1.2600 2.7300 1.6800 2.5500 1.6800 2.5500 2.2100 2.4300 2.2100
                 2.4300 1.5600 2.6100 1.5600 2.6100 0.8150 2.4500 0.8150 2.4500 0.5750 2.5700 0.5750
                 2.5700 0.6950 2.7300 0.6950 2.7300 1.1400 3.1500 1.1400 ;
        POLYGON  2.4900 1.1750 2.3700 1.1750 2.3700 1.0550 1.7700 1.0550 1.7700 1.8150 1.4900 1.8150
                 1.4900 1.9150 1.2500 1.9150 1.2500 1.7950 1.3700 1.7950 1.3700 1.6950 1.6500 1.6950
                 1.6500 1.0550 1.5500 1.0550 1.5500 0.6550 1.3900 0.6550 1.3900 0.4150 1.5100 0.4150
                 1.5100 0.5350 1.6700 0.5350 1.6700 0.9350 2.4900 0.9350 ;
        POLYGON  1.5300 1.5750 1.4100 1.5750 1.4100 1.2950 1.3100 1.2950 1.3100 0.9750 0.2400 0.9750
                 0.2400 1.5550 0.2900 1.5550 0.2900 1.9150 0.1700 1.9150 0.1700 1.6750 0.1200 1.6750
                 0.1200 0.5350 0.3300 0.5350 0.3300 0.4150 0.4500 0.4150 0.4500 0.6550 0.2400 0.6550
                 0.2400 0.8550 1.3100 0.8550 1.3100 0.7750 1.4300 0.7750 1.4300 1.1750 1.5300 1.1750 ;
    END
END MXI2X6

MACRO MXI2X4
    CLASS CORE ;
    FOREIGN MXI2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5950 0.9350 1.7150 1.7550 ;
        RECT  0.9550 1.6350 1.7150 1.7550 ;
        RECT  1.0350 1.5050 1.1550 1.7550 ;
        RECT  0.3900 1.7250 1.0750 1.8450 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.1750 0.8350 1.6050 ;
        RECT  0.6500 1.1750 0.8350 1.5900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0750 1.0500 2.2500 1.4800 ;
        RECT  2.0750 1.0300 2.1950 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6350 0.6800 3.8350 0.8000 ;
        RECT  3.4550 1.3200 3.5750 2.2100 ;
        RECT  2.6250 1.3200 3.5750 1.4400 ;
        RECT  2.6250 1.2300 2.8850 1.4400 ;
        RECT  2.6150 1.4400 2.8750 1.5600 ;
        RECT  2.7550 0.6800 2.8750 1.5600 ;
        RECT  2.6150 1.4400 2.7350 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  4.1950 0.4900 4.4350 0.6100 ;
        RECT  4.3150 -0.1800 4.4350 0.6100 ;
        RECT  3.1150 -0.1800 3.3550 0.3200 ;
        RECT  2.1550 -0.1800 2.2750 0.6700 ;
        RECT  0.6550 -0.1800 0.7750 0.8150 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  3.8750 1.5600 3.9950 2.7900 ;
        RECT  3.0350 1.5600 3.1550 2.7900 ;
        RECT  2.1950 1.6000 2.3150 2.7900 ;
        RECT  0.5550 1.9650 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.7950 0.8600 4.5150 0.8600 4.5150 1.4200 4.4150 1.4200 4.4150 2.2100 4.2950 2.2100
                 4.2950 1.4200 3.6950 1.4200 3.6950 1.3000 4.3950 1.3000 4.3950 0.7400 4.6750 0.7400
                 4.6750 0.6200 4.7950 0.6200 ;
        POLYGON  4.2750 1.1800 4.1550 1.1800 4.1550 0.8500 3.9550 0.8500 3.9550 0.5600 2.5150 0.5600
                 2.5150 0.9100 1.9550 0.9100 1.9550 2.0850 1.3150 2.0850 1.3150 2.2050 1.1950 2.2050
                 1.1950 1.9650 1.8350 1.9650 1.8350 0.8150 1.4550 0.8150 1.4550 0.5750 1.5750 0.5750
                 1.5750 0.6950 1.9550 0.6950 1.9550 0.7900 2.3950 0.7900 2.3950 0.4400 4.0750 0.4400
                 4.0750 0.7300 4.2750 0.7300 ;
        POLYGON  1.4750 1.5150 1.3550 1.5150 1.3550 1.0550 0.2400 1.0550 0.2400 1.8450 0.2550 1.8450
                 0.2550 2.0850 0.1350 2.0850 0.1350 1.9650 0.1200 1.9650 0.1200 0.8150 0.2350 0.8150
                 0.2350 0.5750 0.3550 0.5750 0.3550 0.9350 1.4750 0.9350 ;
    END
END MXI2X4

MACRO MXI2X2
    CLASS CORE ;
    FOREIGN MXI2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 1.3350 1.7400 1.4550 ;
        RECT  1.6200 1.1350 1.7400 1.4550 ;
        RECT  0.9900 1.3350 1.1800 1.5750 ;
        RECT  0.3900 1.5550 1.1100 1.6750 ;
        RECT  0.3900 1.1750 0.5100 1.6750 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6300 1.1750 0.8700 1.4350 ;
        RECT  0.6500 1.1350 0.8700 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1350 2.3200 1.4400 ;
        RECT  2.1000 1.1350 2.2950 1.4600 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6000 1.1750 2.8300 1.4350 ;
        RECT  2.6000 0.8000 2.7200 2.2100 ;
        RECT  2.5500 0.6800 2.6700 0.9200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.0300 -0.1800 3.1500 0.3800 ;
        RECT  2.0700 -0.1800 2.1900 0.7750 ;
        RECT  0.6800 -0.1800 0.8000 0.7750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.0200 1.5600 3.1400 2.7900 ;
        RECT  2.1800 1.5800 2.3000 2.7900 ;
        RECT  0.5800 1.7950 0.7000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.6900 0.8600 3.5700 0.8600 3.5700 1.1950 3.6300 1.1950 3.6300 1.8000 3.5100 1.8000
                 3.5100 1.3150 2.9500 1.3150 2.9500 1.1950 3.4500 1.1950 3.4500 0.7400 3.6900 0.7400 ;
        POLYGON  3.5300 0.5200 3.4100 0.5200 3.4100 0.6200 2.7900 0.6200 2.7900 0.5600 2.4300 0.5600
                 2.4300 1.0150 1.9800 1.0150 1.9800 1.6950 1.4200 1.6950 1.4200 1.8150 1.3500 1.8150
                 1.3500 1.9350 1.2300 1.9350 1.2300 1.6950 1.3000 1.6950 1.3000 1.5750 1.8600 1.5750
                 1.8600 1.0150 1.5950 1.0150 1.5950 0.7750 1.4300 0.7750 1.4300 0.5350 1.5500 0.5350
                 1.5500 0.6550 1.7150 0.6550 1.7150 0.8950 2.3100 0.8950 2.3100 0.4400 2.9100 0.4400
                 2.9100 0.5000 3.2900 0.5000 3.2900 0.4000 3.5300 0.4000 ;
        POLYGON  1.2900 1.1350 1.1700 1.1350 1.1700 1.0150 0.2400 1.0150 0.2400 1.7950 0.2800 1.7950
                 0.2800 2.0350 0.1600 2.0350 0.1600 1.9150 0.1200 1.9150 0.1200 0.7750 0.2600 0.7750
                 0.2600 0.5350 0.3800 0.5350 0.3800 0.8950 1.2900 0.8950 ;
    END
END MXI2X2

MACRO MXI2X1
    CLASS CORE ;
    FOREIGN MXI2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7600 0.5100 1.2100 ;
        RECT  0.3600 0.7600 0.4800 1.3700 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.2300 1.8000 1.4450 ;
        RECT  1.4650 1.2300 1.7250 1.4650 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9900 2.1200 1.1100 ;
        RECT  1.2200 0.9700 2.0150 1.0900 ;
        RECT  1.7550 0.9400 2.0150 1.1100 ;
        RECT  1.4400 0.4100 1.5600 1.0900 ;
        RECT  0.7000 0.4100 1.5600 0.5300 ;
        RECT  0.7000 0.4100 0.8200 1.4300 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 0.6500 1.3200 0.7700 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.9400 0.6500 1.0600 1.6700 ;
        RECT  0.9300 1.5500 1.0500 2.2000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.7800 -0.1800 1.9000 0.8200 ;
        RECT  0.2000 -0.1800 0.3200 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.7100 1.8250 1.8300 2.7900 ;
        RECT  0.2000 1.5500 0.3200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3600 1.8250 2.2500 1.8250 2.2500 2.0650 2.1300 2.0650 2.1300 1.7050 1.2100 1.7050
                 1.2100 1.2300 1.3300 1.2300 1.3300 1.5850 2.2400 1.5850 2.2400 0.8200 2.2000 0.8200
                 2.2000 0.5800 2.3200 0.5800 2.3200 0.7000 2.3600 0.7000 ;
    END
END MXI2X1

MACRO MX4XL
    CLASS CORE ;
    FOREIGN MX4XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7950 1.0400 0.9150 1.4400 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.3200 0.8000 1.7250 ;
        END
    END S1
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0000 1.1600 3.1200 1.6550 ;
        RECT  2.9700 1.1600 3.1200 1.6250 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0750 1.5200 4.3350 1.6700 ;
        RECT  4.0750 1.3300 4.2450 1.6700 ;
        RECT  4.0050 1.3300 4.2450 1.4500 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6000 1.2250 4.7200 1.5150 ;
        RECT  4.3650 1.2250 4.7200 1.4000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5250 0.9700 5.9200 1.1350 ;
        RECT  5.5250 0.9400 5.7850 1.1350 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1050 1.2300 6.3650 1.3800 ;
        RECT  5.4600 1.3300 6.3450 1.4300 ;
        RECT  5.5800 1.3100 6.3650 1.3800 ;
        RECT  5.5800 1.3100 5.7000 2.1700 ;
        RECT  4.1050 2.0500 5.7000 2.1700 ;
        RECT  5.4600 1.3300 5.7000 1.4500 ;
        RECT  3.7650 2.1300 4.2250 2.2500 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.4650 0.2550 1.7050 ;
        RECT  0.1350 0.6800 0.2550 0.9200 ;
        RECT  0.0700 1.4650 0.2200 1.7250 ;
        RECT  0.0950 0.8000 0.2150 1.7250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  5.8400 0.4600 6.0800 0.5800 ;
        RECT  5.9600 -0.1800 6.0800 0.5800 ;
        RECT  4.5400 -0.1800 4.6600 0.8600 ;
        RECT  3.1650 0.6800 3.4050 0.8000 ;
        RECT  3.1650 -0.1800 3.2850 0.8000 ;
        RECT  0.5550 -0.1800 0.6750 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  6.0200 1.7100 6.1400 2.7900 ;
        RECT  4.3450 2.2900 4.5850 2.7900 ;
        RECT  2.8650 2.0200 2.9850 2.7900 ;
        RECT  0.5550 2.0000 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.6050 1.7100 6.5600 1.7100 6.5600 1.8300 6.4400 1.8300 6.4400 1.5900 6.4850 1.5900
                 6.4850 0.8600 6.3800 0.8600 6.3800 0.8200 5.6000 0.8200 5.6000 0.5600 4.9800 0.5600
                 4.9800 1.3100 5.1000 1.3100 5.1000 1.4300 4.8600 1.4300 4.8600 1.1050 4.2200 1.1050
                 4.2200 1.1200 3.8850 1.1200 3.8850 1.3000 3.6000 1.3000 3.6000 1.4200 3.4800 1.4200
                 3.4800 1.1800 3.7650 1.1800 3.7650 0.9850 4.8600 0.9850 4.8600 0.4400 5.2800 0.4400
                 5.2800 0.3600 5.5200 0.3600 5.5200 0.4400 5.7200 0.4400 5.7200 0.7000 6.3800 0.7000
                 6.3800 0.6200 6.5000 0.6200 6.5000 0.7400 6.6050 0.7400 ;
        POLYGON  5.3800 0.8000 5.3400 0.8000 5.3400 1.7100 5.2000 1.7100 5.2000 1.9300 3.9850 1.9300
                 3.9850 2.0100 3.2650 2.0100 3.2650 1.9000 2.4750 1.9000 2.4750 1.3400 2.5350 1.3400
                 2.5350 0.6600 2.6550 0.6600 2.6550 1.4600 2.5950 1.4600 2.5950 1.7800 3.3850 1.7800
                 3.3850 1.8900 3.8650 1.8900 3.8650 1.8100 5.0800 1.8100 5.0800 1.5900 5.2200 1.5900
                 5.2200 0.8000 5.1400 0.8000 5.1400 0.6800 5.3800 0.6800 ;
        POLYGON  4.0200 0.8650 3.6450 0.8650 3.6450 1.0400 3.3600 1.0400 3.3600 1.5400 3.6250 1.5400
                 3.6250 1.6500 3.7450 1.6500 3.7450 1.7700 3.5050 1.7700 3.5050 1.6600 3.2400 1.6600
                 3.2400 1.0400 2.7750 1.0400 2.7750 0.5400 1.8350 0.5400 1.8350 0.6600 1.6950 0.6600
                 1.6950 1.5800 1.7550 1.5800 1.7550 1.7000 1.5150 1.7000 1.5150 1.5800 1.5750 1.5800
                 1.5750 0.5400 1.7150 0.5400 1.7150 0.4200 2.8950 0.4200 2.8950 0.9200 3.5250 0.9200
                 3.5250 0.7450 3.9000 0.7450 3.9000 0.6200 4.0200 0.6200 ;
        POLYGON  2.4150 1.2200 2.3550 1.2200 2.3550 2.1800 1.0350 2.1800 1.0350 0.8000 1.0950 0.8000
                 1.0950 0.6800 1.2150 0.6800 1.2150 0.9200 1.1550 0.9200 1.1550 2.0600 2.2350 2.0600
                 2.2350 0.9800 2.4150 0.9800 ;
        POLYGON  2.1150 1.9400 1.2750 1.9400 1.2750 1.3400 1.3350 1.3400 1.3350 0.5600 0.9150 0.5600
                 0.9150 0.9200 0.5750 0.9200 0.5750 1.2000 0.3350 1.2000 0.3350 1.0800 0.4550 1.0800
                 0.4550 0.8000 0.7950 0.8000 0.7950 0.4400 1.4550 0.4400 1.4550 1.4600 1.3950 1.4600
                 1.3950 1.8200 1.9950 1.8200 1.9950 0.6600 2.1150 0.6600 ;
    END
END MX4XL

MACRO MX4X4
    CLASS CORE ;
    FOREIGN MX4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4550 1.5700 3.6950 1.6900 ;
        RECT  3.4350 0.7400 3.6750 0.8600 ;
        RECT  3.4550 0.7400 3.5750 1.6900 ;
        RECT  2.6800 1.3150 3.5750 1.4350 ;
        RECT  2.5350 1.1750 2.8300 1.3150 ;
        RECT  2.4950 1.5700 2.8000 1.6900 ;
        RECT  2.6800 1.1750 2.8000 1.6900 ;
        RECT  2.5350 0.6800 2.6550 1.3150 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9400 2.0150 1.1550 ;
        RECT  1.7750 0.9400 1.8950 1.3300 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0350 1.0200 4.1550 1.2600 ;
        RECT  3.8400 1.0200 4.1550 1.1450 ;
        RECT  3.8400 0.8850 3.9900 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2350 1.4000 5.4950 1.6700 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8150 1.5200 6.0750 1.6700 ;
        RECT  5.6350 1.5200 6.0750 1.6400 ;
        RECT  5.6350 1.4000 5.7550 1.6400 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2150 1.2300 7.5250 1.4250 ;
        RECT  7.2150 1.2300 7.3350 1.5600 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.2496  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.3867  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9000 1.1750 8.0500 1.4350 ;
        RECT  7.6450 1.1000 8.0200 1.2200 ;
        RECT  7.6450 0.9900 7.7650 1.3400 ;
        RECT  6.7950 0.9900 7.7650 1.1100 ;
        RECT  6.7950 0.9900 6.9150 1.2400 ;
        END
    END S0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.2350 0.7400 7.4750 0.8600 ;
        RECT  7.2350 -0.1800 7.3550 0.8600 ;
        RECT  5.5750 0.6800 5.8150 0.8000 ;
        RECT  5.6950 -0.1800 5.8150 0.8000 ;
        RECT  4.0350 -0.1800 4.1550 0.4000 ;
        RECT  2.9550 -0.1800 3.1950 0.3200 ;
        RECT  1.9950 -0.1800 2.2350 0.3200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.3750 1.9200 7.4950 2.7900 ;
        RECT  5.4350 2.0300 5.6750 2.1500 ;
        RECT  5.4350 2.0300 5.5550 2.7900 ;
        RECT  3.9350 2.0500 4.1750 2.1700 ;
        RECT  3.9350 2.0500 4.0550 2.7900 ;
        RECT  2.9750 2.0500 3.2150 2.1700 ;
        RECT  2.9750 2.0500 3.0950 2.7900 ;
        RECT  2.0150 2.2900 2.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2900 1.9200 7.9150 1.9200 7.9150 2.0400 7.7950 2.0400 7.7950 1.8000 7.0350 1.8000
                 7.0350 2.2200 6.3150 2.2200 6.3150 1.9100 4.9950 1.9100 4.9950 1.6900 4.9350 1.6900
                 4.9350 1.4500 5.0550 1.4500 5.0550 1.5700 5.1150 1.5700 5.1150 1.7900 6.3150 1.7900
                 6.3150 1.0200 6.4350 1.0200 6.4350 2.1000 6.9150 2.1000 6.9150 1.6600 6.8150 1.6600
                 6.8150 1.5400 7.0550 1.5400 7.0550 1.6800 8.1700 1.6800 8.1700 0.8600 7.6550 0.8600
                 7.6550 0.7400 8.2900 0.7400 ;
        POLYGON  6.7950 1.9800 6.5550 1.9800 6.5550 0.9000 6.1450 0.9000 6.1450 1.0400 5.2300 1.0400
                 5.2300 0.5600 4.3950 0.5600 4.3950 0.6400 3.7950 0.6400 3.7950 0.6200 3.0000 0.6200
                 3.0000 0.5600 1.7550 0.5600 1.7550 0.4800 1.2150 0.4800 1.2150 0.6000 1.2850 0.6000
                 1.2850 1.5600 1.3850 1.5600 1.3850 1.6900 1.1450 1.6900 1.1450 1.5600 1.1650 1.5600
                 1.1650 0.7200 1.0950 0.7200 1.0950 0.3600 1.8750 0.3600 1.8750 0.4400 3.1200 0.4400
                 3.1200 0.5000 3.9150 0.5000 3.9150 0.5200 4.2750 0.5200 4.2750 0.4400 5.3500 0.4400
                 5.3500 0.9200 6.0250 0.9200 6.0250 0.7800 6.5550 0.7800 6.5550 0.6800 6.6750 0.6800
                 6.6750 1.8600 6.7950 1.8600 ;
        POLYGON  6.1550 1.4000 5.9150 1.4000 5.9150 1.2800 4.6350 1.2800 4.6350 1.4800 4.5150 1.4800
                 4.5150 1.1600 6.1550 1.1600 ;
        POLYGON  5.0550 0.9200 4.3950 0.9200 4.3950 1.8100 4.8750 1.8100 4.8750 1.9800 4.6350 1.9800
                 4.6350 1.9300 2.4700 1.9300 2.4700 2.1700 1.4100 2.1700 1.4100 2.2500 0.3650 2.2500
                 0.3650 1.4000 0.1050 1.4000 0.1050 0.6800 0.1350 0.6800 0.1350 0.5600 0.2550 0.5600
                 0.2550 0.8000 0.2250 0.8000 0.2250 1.2800 0.4850 1.2800 0.4850 2.1300 1.2900 2.1300
                 1.2900 2.0500 2.3500 2.0500 2.3500 1.8100 4.2750 1.8100 4.2750 0.8000 4.9350 0.8000
                 4.9350 0.6800 5.0550 0.6800 ;
        POLYGON  2.4150 1.4500 2.3750 1.4500 2.3750 1.5700 2.2300 1.5700 2.2300 1.9300 0.9050 1.9300
                 0.9050 2.0100 0.7850 2.0100 0.7850 1.6200 0.6150 1.6200 0.6150 0.6000 0.7350 0.6000
                 0.7350 1.5000 0.9050 1.5000 0.9050 1.8100 2.1100 1.8100 2.1100 1.4500 2.2550 1.4500
                 2.2550 1.3300 2.2950 1.3300 2.2950 1.1700 2.4150 1.1700 ;
        POLYGON  1.7750 1.6900 1.5150 1.6900 1.5150 1.4000 1.4050 1.4000 1.4050 1.1600 1.5150 1.1600
                 1.5150 0.6000 1.6350 0.6000 1.6350 1.5700 1.7750 1.5700 ;
        POLYGON  1.0450 1.3800 0.9250 1.3800 0.9250 1.2600 0.8550 1.2600 0.8550 0.4800 0.4950 0.4800
                 0.4950 1.1600 0.3450 1.1600 0.3450 0.9200 0.3750 0.9200 0.3750 0.3600 0.9750 0.3600
                 0.9750 1.1400 1.0450 1.1400 ;
    END
END MX4X4

MACRO MX4X2
    CLASS CORE ;
    FOREIGN MX4X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.2500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7900 0.8850 1.9600 1.1550 ;
        RECT  1.7300 1.0350 1.8700 1.2850 ;
        END
    END S1
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9500 1.0800 3.0700 1.3200 ;
        RECT  2.6800 1.1750 3.0700 1.2950 ;
        RECT  2.6800 1.1750 2.8300 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1300 1.4000 4.3000 1.8350 ;
        RECT  4.1700 1.3800 4.3000 1.8350 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4900 1.3800 4.6700 1.6300 ;
        RECT  4.4200 1.4600 4.6250 1.7250 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0500 1.2000 6.3650 1.4150 ;
        RECT  6.0500 1.2000 6.1700 1.5600 ;
        END
    END D
    PIN S0
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.2976  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.6533  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4850 1.1750 6.8900 1.4350 ;
        RECT  6.4850 0.9600 6.6050 1.4350 ;
        RECT  5.7100 0.9600 6.6050 1.0800 ;
        RECT  5.7100 0.9600 5.8300 1.2200 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3500 1.5700 2.5900 1.6900 ;
        RECT  2.4700 0.6600 2.5900 1.0250 ;
        RECT  2.4200 0.8850 2.5400 1.6900 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.2500 0.1800 ;
        RECT  6.1500 0.7200 6.3900 0.8400 ;
        RECT  6.1500 -0.1800 6.2700 0.8400 ;
        RECT  4.4500 0.5400 4.6900 0.6600 ;
        RECT  4.5700 -0.1800 4.6900 0.6600 ;
        RECT  2.9500 -0.1800 3.0700 0.3800 ;
        RECT  1.9900 -0.1800 2.1100 0.5250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.2500 2.7900 ;
        RECT  6.2100 1.9200 6.3300 2.7900 ;
        RECT  4.3400 2.1950 4.5800 2.7900 ;
        RECT  2.8300 2.0500 3.0700 2.1700 ;
        RECT  2.8300 2.0500 2.9500 2.7900 ;
        RECT  1.8700 2.2900 2.1100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.1300 1.9200 6.7500 1.9200 6.7500 2.0400 6.6300 2.0400 6.6300 1.8000 5.9100 1.8000
                 5.9100 2.2200 5.1900 2.2200 5.1900 2.0750 3.8900 2.0750 3.8900 1.7400 3.8400 1.7400
                 3.8400 1.4800 3.9600 1.4800 3.9600 1.6200 4.0100 1.6200 4.0100 1.9550 5.1900 1.9550
                 5.1900 1.0000 5.3100 1.0000 5.3100 2.1000 5.7900 2.1000 5.7900 1.7400 5.7300 1.7400
                 5.7300 1.4600 5.8500 1.4600 5.8500 1.6200 5.9100 1.6200 5.9100 1.6800 7.0100 1.6800
                 7.0100 1.0550 6.7250 1.0550 6.7250 0.6600 6.8450 0.6600 6.8450 0.9350 7.1300 0.9350 ;
        POLYGON  5.6700 1.9800 5.4300 1.9800 5.4300 0.8800 4.9650 0.8800 4.9650 0.9000 4.0500 0.9000
                 4.0500 0.5400 3.3750 0.5400 3.3750 0.6200 2.7100 0.6200 2.7100 0.5400 2.3500 0.5400
                 2.3500 0.7650 1.7500 0.7650 1.7500 0.4900 1.2150 0.4900 1.2150 0.9300 1.2400 0.9300
                 1.2400 1.6500 1.1800 1.6500 1.1800 1.7700 1.0600 1.7700 1.0600 1.5300 1.1200 1.5300
                 1.1200 1.0500 1.0950 1.0500 1.0950 0.3700 1.8700 0.3700 1.8700 0.6450 2.2300 0.6450
                 2.2300 0.4200 2.8300 0.4200 2.8300 0.5000 3.2550 0.5000 3.2550 0.4200 4.1700 0.4200
                 4.1700 0.7800 4.8450 0.7800 4.8450 0.7600 5.4300 0.7600 5.4300 0.6600 5.5500 0.6600
                 5.5500 1.8600 5.6700 1.8600 ;
        POLYGON  5.0300 1.4200 4.7900 1.4200 4.7900 1.2600 3.7200 1.2600 3.7200 1.5800 3.5500 1.5800
                 3.5500 1.7000 3.4300 1.7000 3.4300 1.4600 3.6000 1.4600 3.6000 1.1400 3.9700 1.1400
                 3.9700 1.0200 4.0900 1.0200 4.0900 1.1400 5.0300 1.1400 ;
        POLYGON  3.9300 0.9000 3.4800 0.9000 3.4800 1.3400 3.3100 1.3400 3.3100 1.8200 3.6500 1.8200
                 3.6500 1.8600 3.7700 1.8600 3.7700 1.9800 3.5300 1.9800 3.5300 1.9400 3.1900 1.9400
                 3.1900 1.9300 2.2500 1.9300 2.2500 2.1700 1.6650 2.1700 1.6650 2.2500 0.2200 2.2500
                 0.2200 1.4400 0.0800 1.4400 0.0800 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000
                 0.2550 0.8400 0.2000 0.8400 0.2000 1.3200 0.3400 1.3200 0.3400 2.1300 1.5450 2.1300
                 1.5450 2.0500 2.1300 2.0500 2.1300 1.8100 3.1900 1.8100 3.1900 1.2200 3.3600 1.2200
                 3.3600 0.7800 3.8100 0.7800 3.8100 0.6600 3.9300 0.6600 ;
        POLYGON  2.2700 1.4100 2.2300 1.4100 2.2300 1.5300 2.0100 1.5300 2.0100 1.9300 1.4250 1.9300
                 1.4250 2.0100 0.6400 2.0100 0.6400 1.6400 0.6150 1.6400 0.6150 0.6000 0.7350 0.6000
                 0.7350 1.5200 0.7600 1.5200 0.7600 1.8900 1.3050 1.8900 1.3050 1.8100 1.8900 1.8100
                 1.8900 1.4100 2.1100 1.4100 2.1100 1.2900 2.1500 1.2900 2.1500 1.1700 2.2700 1.1700 ;
        POLYGON  1.6300 0.9150 1.5100 0.9150 1.5100 1.5700 1.6300 1.5700 1.6300 1.6900 1.3900 1.6900
                 1.3900 1.4100 1.3600 1.4100 1.3600 1.1700 1.3900 1.1700 1.3900 0.7950 1.5100 0.7950
                 1.5100 0.6100 1.6300 0.6100 ;
        POLYGON  1.0000 1.4100 0.8800 1.4100 0.8800 1.2900 0.8550 1.2900 0.8550 0.4800 0.4950 0.4800
                 0.4950 1.2000 0.3200 1.2000 0.3200 0.9600 0.3750 0.9600 0.3750 0.3600 0.9750 0.3600
                 0.9750 1.1700 1.0000 1.1700 ;
    END
END MX4X2

MACRO MX4X1
    CLASS CORE ;
    FOREIGN MX4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.2500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9450 1.0050 1.1850 1.2200 ;
        RECT  0.8850 0.9400 1.1450 1.1800 ;
        END
    END S1
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3450 1.2600 3.5850 1.4500 ;
        RECT  3.2050 1.1650 3.4650 1.3800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7050 1.2700 4.8250 1.5400 ;
        RECT  4.5050 1.4200 4.8250 1.5400 ;
        RECT  4.3650 1.5200 4.6250 1.6700 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 1.5200 5.2050 1.6700 ;
        RECT  5.0650 1.2500 5.1850 1.6700 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.2450 1.0050 6.5050 1.1600 ;
        RECT  6.1050 0.9400 6.3650 1.1250 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6850 1.2300 6.9450 1.3800 ;
        RECT  5.9250 1.3100 6.8250 1.4300 ;
        RECT  6.0450 1.3100 6.1650 2.1700 ;
        RECT  4.6050 2.0500 6.1650 2.1700 ;
        RECT  4.2450 2.1300 4.7250 2.2500 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3650 1.3400 0.4850 1.9900 ;
        RECT  0.2900 0.5900 0.4100 1.4600 ;
        RECT  0.0700 0.8850 0.4100 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.2500 0.1800 ;
        RECT  6.3050 0.4600 6.5450 0.5800 ;
        RECT  6.4250 -0.1800 6.5450 0.5800 ;
        RECT  5.0050 -0.1800 5.1250 0.8600 ;
        RECT  3.6050 0.5300 3.8450 0.6500 ;
        RECT  3.6050 -0.1800 3.7250 0.6500 ;
        RECT  0.6500 0.4600 0.8900 0.5800 ;
        RECT  0.6500 -0.1800 0.7700 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.2500 2.7900 ;
        RECT  6.4850 1.7100 6.6050 2.7900 ;
        RECT  4.8450 2.2900 5.0850 2.7900 ;
        RECT  3.3650 2.0200 3.4850 2.7900 ;
        RECT  0.7850 1.3400 0.9050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.1850 1.6700 7.0250 1.6700 7.0250 1.8300 6.9050 1.8300 6.9050 1.5500 7.0650 1.5500
                 7.0650 0.8600 6.8450 0.8600 6.8450 0.8200 6.0650 0.8200 6.0650 0.5600 5.4450 0.5600
                 5.4450 1.3100 5.5650 1.3100 5.5650 1.4300 5.3250 1.4300 5.3250 1.1300 4.5850 1.1300
                 4.5850 1.3000 4.0650 1.3000 4.0650 1.4200 3.9450 1.4200 3.9450 1.1800 4.4450 1.1800
                 4.4450 1.0100 5.3250 1.0100 5.3250 0.4400 5.7450 0.4400 5.7450 0.3600 5.9850 0.3600
                 5.9850 0.4400 6.1850 0.4400 6.1850 0.7000 6.8450 0.7000 6.8450 0.6200 6.9650 0.6200
                 6.9650 0.7400 7.1850 0.7400 ;
        POLYGON  5.8450 0.8000 5.8050 0.8000 5.8050 1.9300 4.4850 1.9300 4.4850 2.0100 3.6050 2.0100
                 3.6050 1.9000 2.8100 1.9000 2.8100 1.2200 2.9300 1.2200 2.9300 0.8600 2.8100 0.8600
                 2.8100 0.6000 2.9300 0.6000 2.9300 0.7400 3.0500 0.7400 3.0500 1.3400 2.9300 1.3400
                 2.9300 1.7800 3.7250 1.7800 3.7250 1.8900 4.3650 1.8900 4.3650 1.8100 5.6850 1.8100
                 5.6850 0.8000 5.6050 0.8000 5.6050 0.6800 5.8450 0.6800 ;
        POLYGON  4.4850 0.8900 3.8250 0.8900 3.8250 1.5400 4.1250 1.5400 4.1250 1.6500 4.2450 1.6500
                 4.2450 1.7700 4.0050 1.7700 4.0050 1.6600 3.7050 1.6600 3.7050 0.8900 3.3650 0.8900
                 3.3650 0.4800 2.0900 0.4800 2.0900 1.6400 1.8500 1.6400 1.8500 1.5200 1.9700 1.5200
                 1.9700 0.3600 3.4850 0.3600 3.4850 0.7700 4.3650 0.7700 4.3650 0.6200 4.4850 0.6200 ;
        POLYGON  2.8100 1.1000 2.6900 1.1000 2.6900 2.1200 1.2650 2.1200 1.2650 1.4600 1.3050 1.4600
                 1.3050 0.7700 1.2500 0.7700 1.2500 0.6500 1.4900 0.6500 1.4900 0.7700 1.4250 0.7700
                 1.4250 1.5800 1.3850 1.5800 1.3850 2.0000 2.5700 2.0000 2.5700 0.9800 2.8100 0.9800 ;
        POLYGON  2.5100 0.8400 2.4500 0.8400 2.4500 1.8800 1.6100 1.8800 1.6100 0.5300 1.1300 0.5300
                 1.1300 0.8200 0.7650 0.8200 0.7650 1.1500 0.6450 1.1500 0.6450 0.7000 1.0100 0.7000
                 1.0100 0.4100 1.7300 0.4100 1.7300 1.7600 2.3300 1.7600 2.3300 0.7200 2.3900 0.7200
                 2.3900 0.6000 2.5100 0.6000 ;
    END
END MX4X1

MACRO MX3XL
    CLASS CORE ;
    FOREIGN MX3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7100 1.2500 0.8300 1.5550 ;
        RECT  0.6500 1.4350 0.8000 1.7500 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.7850 2.5400 1.1800 ;
        RECT  2.3800 1.0600 2.5000 1.4700 ;
        END
    END S1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7200 0.7850 2.8400 1.2700 ;
        RECT  2.6800 0.7700 2.8300 1.2300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8000 1.0100 4.0400 1.1300 ;
        RECT  3.8400 1.0100 3.9900 1.4350 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1300 1.4650 4.2800 1.7250 ;
        RECT  4.1400 1.4350 4.2600 1.7250 ;
        RECT  3.5600 1.5550 4.2800 1.6750 ;
        RECT  3.5600 1.2500 3.6800 1.6750 ;
        RECT  3.4800 1.1100 3.6000 1.3700 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 1.8500 0.4100 1.9700 ;
        RECT  0.2900 0.6100 0.4100 1.9700 ;
        RECT  0.0700 0.8850 0.4100 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  3.9800 -0.1800 4.1000 0.6500 ;
        RECT  2.7000 -0.1800 2.8200 0.6500 ;
        RECT  0.7100 -0.1800 0.8300 0.8500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  3.9800 1.9700 4.1000 2.7900 ;
        RECT  2.7000 1.9700 2.8200 2.7900 ;
        RECT  0.6500 1.9100 0.7700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.5200 2.0900 4.4000 2.0900 4.4000 0.8900 3.6800 0.8900 3.6800 0.9900 3.3600 0.9900
                 3.3600 1.4900 3.4400 1.4900 3.4400 1.6100 3.2000 1.6100 3.2000 1.4900 3.2400 1.4900
                 3.2400 0.8700 3.4400 0.8700 3.4400 0.8100 3.5600 0.8100 3.5600 0.7700 4.4000 0.7700
                 4.4000 0.4100 4.5200 0.4100 ;
        POLYGON  3.4600 0.6500 3.3200 0.6500 3.3200 0.7500 3.0800 0.7500 3.0800 1.7300 3.4400 1.7300
                 3.4400 1.8500 3.4600 1.8500 3.4600 2.0900 3.3400 2.0900 3.3400 1.9700 3.3200 1.9700
                 3.3200 1.8500 2.0900 1.8500 2.0900 1.9700 1.8300 1.9700 1.8300 1.8500 1.9700 1.8500
                 1.9700 0.8500 1.8900 0.8500 1.8900 0.6100 2.0100 0.6100 2.0100 0.7300 2.0900 0.7300
                 2.0900 1.7300 2.9600 1.7300 2.9600 0.6300 3.2000 0.6300 3.2000 0.5300 3.3400 0.5300
                 3.3400 0.4100 3.4600 0.4100 ;
        POLYGON  2.4000 0.6500 2.2800 0.6500 2.2800 0.4900 1.7700 0.4900 1.7700 0.9700 1.8500 0.9700
                 1.8500 1.2100 1.7700 1.2100 1.7700 1.5700 1.7100 1.5700 1.7100 2.0900 2.2800 2.0900
                 2.2800 1.9700 2.4000 1.9700 2.4000 2.2100 1.5900 2.2100 1.5900 1.5700 1.3100 1.5700
                 1.3100 1.6900 1.1900 1.6900 1.1900 1.4500 1.6500 1.4500 1.6500 0.3700 2.4000 0.3700 ;
        POLYGON  1.5300 1.1100 1.0700 1.1100 1.0700 1.8100 1.3500 1.8100 1.3500 1.8500 1.4700 1.8500
                 1.4700 1.9700 1.2300 1.9700 1.2300 1.9300 0.9500 1.9300 0.9500 1.1100 0.5300 1.1100
                 0.5300 0.9900 1.4100 0.9900 1.4100 0.6100 1.5300 0.6100 ;
    END
END MX3XL

MACRO MX3X4
    CLASS CORE ;
    FOREIGN MX3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.0400 2.3500 1.2450 ;
        RECT  2.1000 1.0400 2.2500 1.4350 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8400 0.7600 3.9900 1.1450 ;
        RECT  3.8200 1.0250 3.9400 1.4200 ;
        END
    END S1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1600 0.7900 4.2800 1.3200 ;
        RECT  4.1300 0.7900 4.2800 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2800 1.1450 5.5200 1.3450 ;
        RECT  5.2900 1.0700 5.4400 1.4600 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 1.5800 5.7800 1.7000 ;
        RECT  5.6600 1.4400 5.7800 1.7000 ;
        RECT  5.5800 1.4650 5.7300 1.7250 ;
        RECT  5.0000 1.4600 5.1200 1.7000 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6700 1.2800 1.7900 2.1700 ;
        RECT  1.5000 0.5600 1.7900 0.6800 ;
        RECT  1.6700 0.4400 1.7900 0.6800 ;
        RECT  0.6500 1.2800 1.7900 1.4000 ;
        RECT  0.8300 0.7700 1.6200 0.8900 ;
        RECT  1.5000 0.5600 1.6200 0.8900 ;
        RECT  0.8300 0.6000 0.9500 2.1700 ;
        RECT  0.6500 1.1750 0.9500 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.5000 -0.1800 5.6200 0.6400 ;
        RECT  4.2200 -0.1800 4.3400 0.6400 ;
        RECT  2.0900 -0.1800 2.2100 0.6500 ;
        RECT  1.2500 -0.1800 1.3700 0.6500 ;
        RECT  0.4100 -0.1800 0.5300 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.4400 1.9600 5.6800 2.0800 ;
        RECT  5.4400 1.9600 5.5600 2.7900 ;
        RECT  4.0800 1.9000 4.2000 2.7900 ;
        RECT  2.0900 1.5550 2.2100 2.7900 ;
        RECT  1.2500 1.5200 1.3700 2.7900 ;
        RECT  0.4100 1.5200 0.5300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.1000 1.9600 5.8600 1.9600 5.8600 1.8400 5.9000 1.8400 5.9000 0.9500 5.1200 0.9500
                 5.1200 1.3400 4.7600 1.3400 4.7600 1.5400 4.6400 1.5400 4.6400 1.2200 5.0000 1.2200
                 5.0000 0.7600 5.1200 0.7600 5.1200 0.8300 5.9000 0.8300 5.9000 0.5200 5.9200 0.5200
                 5.9200 0.4000 6.0400 0.4000 6.0400 0.6400 6.0200 0.6400 6.0200 1.8400 6.1000 1.8400 ;
        POLYGON  4.9800 0.6400 4.8800 0.6400 4.8800 1.1000 4.5200 1.1000 4.5200 1.6600 4.7800 1.6600
                 4.7800 1.8400 4.9000 1.8400 4.9000 1.9600 4.6600 1.9600 4.6600 1.7800 3.4500 1.7800
                 3.4500 2.0100 3.2100 2.0100 3.2100 1.5800 3.4900 1.5800 3.4900 0.8400 3.4100 0.8400
                 3.4100 0.6000 3.5300 0.6000 3.5300 0.7200 3.6100 0.7200 3.6100 1.6600 4.4000 1.6600
                 4.4000 0.9800 4.7600 0.9800 4.7600 0.5200 4.8600 0.5200 4.8600 0.4000 4.9800 0.4000 ;
        POLYGON  3.9200 0.6400 3.8000 0.6400 3.8000 0.4800 3.2900 0.4800 3.2900 0.9600 3.3700 0.9600
                 3.3700 1.2000 3.2900 1.2000 3.2900 1.4600 3.0900 1.4600 3.0900 2.1300 3.6000 2.1300
                 3.6000 1.9600 3.8400 1.9600 3.8400 2.0800 3.7200 2.0800 3.7200 2.2500 2.9700 2.2500
                 2.9700 1.4000 2.7100 1.4000 2.7100 1.1600 2.8300 1.1600 2.8300 1.2800 3.1700 1.2800
                 3.1700 0.3600 3.9200 0.3600 ;
        POLYGON  3.0500 0.9200 2.5900 0.9200 2.5900 1.5200 2.8500 1.5200 2.8500 2.1700 2.7300 2.1700
                 2.7300 1.6400 2.4700 1.6400 2.4700 0.9200 1.9800 0.9200 1.9800 1.1000 1.7400 1.1000
                 1.7400 0.8000 2.9300 0.8000 2.9300 0.6000 3.0500 0.6000 ;
    END
END MX3X4

MACRO MX3X2
    CLASS CORE ;
    FOREIGN MX3X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2300 1.2650 1.3900 ;
        RECT  1.1450 1.1300 1.2650 1.3900 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7100 0.7600 2.8300 1.4300 ;
        RECT  2.6800 0.7600 2.8300 1.1600 ;
        END
    END S1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.8850 3.3150 1.0600 ;
        RECT  3.1950 0.8200 3.3150 1.0600 ;
        RECT  2.9700 0.8850 3.1200 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4200 1.0850 4.5700 1.4600 ;
        RECT  4.2950 1.1100 4.5700 1.3000 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7100 1.4650 4.8600 1.7250 ;
        RECT  4.7100 1.4600 4.8300 1.7250 ;
        RECT  4.0150 1.5800 4.8600 1.7000 ;
        RECT  4.0150 1.4600 4.1350 1.7000 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6450 1.3500 0.7650 2.1600 ;
        RECT  0.4850 0.6500 0.7650 0.7700 ;
        RECT  0.6450 0.5300 0.7650 0.7700 ;
        RECT  0.4850 1.3500 0.7650 1.4700 ;
        RECT  0.3050 1.2300 0.6050 1.3800 ;
        RECT  0.4850 0.6500 0.6050 1.4700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  4.4150 -0.1800 4.5350 0.6400 ;
        RECT  3.1350 -0.1800 3.2550 0.6400 ;
        RECT  1.0050 0.4800 1.2450 0.6000 ;
        RECT  1.0050 -0.1800 1.1250 0.6000 ;
        RECT  0.2250 -0.1800 0.3450 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  4.5150 1.9400 4.6350 2.7900 ;
        RECT  3.1950 1.9400 3.3150 2.7900 ;
        RECT  1.0650 1.5100 1.1850 2.7900 ;
        RECT  0.2250 1.5100 0.3450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.1000 1.9650 5.0550 1.9650 5.0550 2.0850 4.9350 2.0850 4.9350 1.8450 4.9800 1.8450
                 4.9800 0.9650 4.0550 0.9650 4.0550 1.0000 3.8950 1.0000 3.8950 1.4600 3.7950 1.4600
                 3.7950 1.5800 3.6750 1.5800 3.6750 1.3400 3.7750 1.3400 3.7750 0.8450 3.9350 0.8450
                 3.9350 0.7600 4.0550 0.7600 4.0550 0.8450 4.9800 0.8450 4.9800 0.6400 4.8350 0.6400
                 4.8350 0.4000 4.9550 0.4000 4.9550 0.5200 5.1000 0.5200 ;
        POLYGON  3.9550 2.0600 3.8350 2.0600 3.8350 1.9400 3.7750 1.9400 3.7750 1.8200 2.4050 1.8200
                 2.4050 1.6900 2.1850 1.6900 2.1850 1.5700 2.4050 1.5700 2.4050 0.7900 2.2650 0.7900
                 2.2650 0.6700 2.5250 0.6700 2.5250 1.7000 3.4350 1.7000 3.4350 1.1000 3.5350 1.1000
                 3.5350 0.5200 3.7750 0.5200 3.7750 0.4000 3.8950 0.4000 3.8950 0.6400 3.6550 0.6400
                 3.6550 1.2200 3.5550 1.2200 3.5550 1.7000 3.8950 1.7000 3.8950 1.8200 3.9550 1.8200 ;
        POLYGON  2.9550 2.0600 1.9450 2.0600 1.9450 1.2900 1.7450 1.2900 1.7450 1.4100 1.6250 1.4100
                 1.6250 1.1700 2.1650 1.1700 2.1650 1.0300 2.0250 1.0300 2.0250 0.4300 2.7150 0.4300
                 2.7150 0.4000 2.8350 0.4000 2.8350 0.6400 2.7150 0.6400 2.7150 0.5500 2.1450 0.5500
                 2.1450 0.9100 2.2850 0.9100 2.2850 1.4500 2.0650 1.4500 2.0650 1.9400 2.9550 1.9400 ;
        POLYGON  1.9050 1.0100 1.5050 1.0100 1.5050 1.5300 1.8250 1.5300 1.8250 1.7700 1.7050 1.7700
                 1.7050 1.6500 1.3850 1.6500 1.3850 1.0100 0.9650 1.0100 0.9650 1.1100 0.7250 1.1100
                 0.7250 0.8900 1.7850 0.8900 1.7850 0.6100 1.9050 0.6100 ;
    END
END MX3X2

MACRO MX3X1
    CLASS CORE ;
    FOREIGN MX3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8200 1.1900 1.0900 1.4500 ;
        RECT  0.9400 1.1750 1.0900 1.4500 ;
        END
    END C
    PIN S1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 0.8850 2.2500 1.3550 ;
        RECT  2.1300 0.8550 2.2500 1.3550 ;
        END
    END S1
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6950 1.0400 2.8150 1.2800 ;
        RECT  2.4200 1.0400 2.8150 1.1600 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8200 1.1100 4.0600 1.3000 ;
        RECT  3.8400 1.0800 3.9900 1.4550 ;
        END
    END A
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2200 1.5200 4.6250 1.6700 ;
        RECT  4.2200 1.5000 4.4600 1.6700 ;
        RECT  3.5400 1.5750 4.3400 1.6950 ;
        RECT  3.5400 1.4600 3.6600 1.7000 ;
        END
    END S0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2000 1.3000 0.3200 2.2100 ;
        RECT  0.2000 0.6800 0.3200 0.9400 ;
        RECT  0.1600 0.8200 0.2800 1.4200 ;
        RECT  0.0700 0.8850 0.2800 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  4.1950 0.5200 4.4350 0.6400 ;
        RECT  4.1950 -0.1800 4.3150 0.6400 ;
        RECT  2.9750 -0.1800 3.0950 0.7000 ;
        RECT  0.5600 0.5500 0.8000 0.6700 ;
        RECT  0.5600 -0.1800 0.6800 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  4.0400 1.9000 4.1600 2.7900 ;
        RECT  2.7600 1.9000 2.8800 2.7900 ;
        RECT  0.6200 1.7200 0.7400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8650 1.9100 4.5800 1.9100 4.5800 2.0300 4.4600 2.0300 4.4600 1.7900 4.7450 1.7900
                 4.7450 0.9600 3.7000 0.9600 3.7000 1.3400 3.2950 1.3400 3.2950 1.4800 3.1750 1.4800
                 3.1750 1.2200 3.5800 1.2200 3.5800 0.8400 4.7450 0.8400 4.7450 0.7000 4.6750 0.7000
                 4.6750 0.4600 4.7950 0.4600 4.7950 0.5800 4.8650 0.5800 ;
        POLYGON  3.7950 0.6400 3.4600 0.6400 3.4600 1.1000 3.0550 1.1000 3.0550 1.6600 3.4200 1.6600
                 3.4200 1.8200 3.5200 1.8200 3.5200 2.0600 3.4000 2.0600 3.4000 1.9400 3.3000 1.9400
                 3.3000 1.7800 2.1300 1.7800 2.1300 1.9000 1.8600 1.9000 1.8600 0.6000 2.1000 0.6000
                 2.1000 0.7200 1.9800 0.7200 1.9800 1.6600 2.9350 1.6600 2.9350 0.9800 3.3400 0.9800
                 3.3400 0.5200 3.7950 0.5200 ;
        POLYGON  2.6750 0.7000 2.5550 0.7000 2.5550 0.4800 1.7400 0.4800 1.7400 2.0200 2.3400 2.0200
                 2.3400 1.9000 2.4600 1.9000 2.4600 2.1400 1.6200 2.1400 1.6200 1.6400 1.4500 1.6400
                 1.4500 1.4000 1.6200 1.4000 1.6200 1.0400 1.5000 1.0400 1.5000 0.9200 1.6200 0.9200
                 1.6200 0.3600 2.6750 0.3600 ;
        POLYGON  1.5000 0.7200 1.3800 0.7200 1.3800 1.0550 1.3300 1.0550 1.3300 1.7800 1.5000 1.7800
                 1.5000 1.9000 1.2100 1.9000 1.2100 1.0550 0.7000 1.0550 0.7000 1.1800 0.4000 1.1800
                 0.4000 1.0600 0.5800 1.0600 0.5800 0.9350 1.2600 0.9350 1.2600 0.6000 1.5000 0.6000 ;
    END
END MX3X1

MACRO MX2XL
    CLASS CORE ;
    FOREIGN MX2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9700 1.2550 1.2500 1.3750 ;
        RECT  0.4100 1.6950 1.0900 1.8150 ;
        RECT  0.9700 1.2550 1.0900 1.8150 ;
        RECT  0.3600 1.4750 0.5300 1.7250 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1050 0.8500 1.5750 ;
        RECT  0.7300 1.0750 0.8500 1.5750 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9100 1.3150 2.2500 1.4350 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.9100 1.3150 2.0300 1.5550 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.1750 2.5400 1.4350 ;
        RECT  2.4100 1.1750 2.5300 2.0550 ;
        RECT  2.3700 0.4750 2.4900 1.3150 ;
        RECT  2.3900 1.1750 2.5300 1.5550 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.8900 0.5350 2.1300 0.6550 ;
        RECT  1.8900 -0.1800 2.0100 0.6550 ;
        RECT  0.6700 -0.1800 0.7900 0.7150 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.9900 1.9350 2.1100 2.7900 ;
        RECT  0.7100 1.9350 0.8300 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2500 1.0550 1.7900 1.0550 1.7900 1.9750 1.5300 1.9750 1.5300 1.9950 1.2900 1.9950
                 1.2900 1.8750 1.4100 1.8750 1.4100 1.8550 1.6700 1.8550 1.6700 1.0550 1.6100 1.0550
                 1.6100 0.7150 1.3100 0.7150 1.3100 0.4750 1.4300 0.4750 1.4300 0.5950 1.7300 0.5950
                 1.7300 0.9350 2.1300 0.9350 2.1300 0.8150 2.2500 0.8150 ;
        POLYGON  1.5500 1.7350 1.4300 1.7350 1.4300 1.2950 1.3700 1.2950 1.3700 1.0750 1.1500 1.0750
                 1.1500 0.9550 0.2400 0.9550 0.2400 1.9350 0.4100 1.9350 0.4100 2.1750 0.2900 2.1750
                 0.2900 2.0550 0.1200 2.0550 0.1200 0.5950 0.2500 0.5950 0.2500 0.4750 0.3700 0.4750
                 0.3700 0.7150 0.2400 0.7150 0.2400 0.8350 1.4900 0.8350 1.4900 1.1750 1.5500 1.1750 ;
    END
END MX2XL

MACRO MX2X8
    CLASS CORE ;
    FOREIGN MX2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.8000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 1.1200 1.5050 1.2400 ;
        RECT  0.6450 1.5000 1.3850 1.6200 ;
        RECT  1.2650 1.1200 1.3850 1.6200 ;
        RECT  0.6450 1.1750 0.7650 1.6200 ;
        RECT  0.3600 1.1750 0.7650 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1100 1.1450 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0800 2.5400 1.4600 ;
        RECT  2.2800 1.0800 2.5400 1.2750 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7250 0.7650 5.4650 0.8850 ;
        RECT  5.3450 0.6450 5.4650 0.8850 ;
        RECT  5.3400 0.7650 5.4600 2.2050 ;
        RECT  2.9700 1.2250 5.4600 1.3450 ;
        RECT  4.4450 0.7150 4.6850 0.8850 ;
        RECT  4.5000 1.2250 4.6200 2.2050 ;
        RECT  3.6050 0.7150 3.8450 0.8350 ;
        RECT  3.6600 1.2250 3.7800 2.2100 ;
        RECT  2.9700 1.1750 3.1200 1.4350 ;
        RECT  2.8200 1.3450 3.0900 1.4650 ;
        RECT  2.9700 0.6000 3.0900 1.4650 ;
        RECT  2.7650 0.6000 3.0900 0.7200 ;
        RECT  2.8200 1.3450 2.9400 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.8000 0.1800 ;
        RECT  4.9250 -0.1800 5.0450 0.6450 ;
        RECT  4.0850 -0.1800 4.2050 0.6450 ;
        RECT  3.2450 -0.1800 3.3650 0.6450 ;
        RECT  2.3450 0.4600 2.5850 0.5800 ;
        RECT  2.3450 -0.1800 2.4650 0.5800 ;
        RECT  0.8250 -0.1800 0.9450 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.8000 2.7900 ;
        RECT  4.9200 1.4650 5.0400 2.7900 ;
        RECT  4.0800 1.4650 4.2000 2.7900 ;
        RECT  3.2400 1.4650 3.3600 2.7900 ;
        RECT  2.4000 1.5800 2.5200 2.7900 ;
        RECT  0.9600 1.7400 1.2000 2.1400 ;
        RECT  0.9600 1.7400 1.0800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.8000 1.2150 2.6800 1.2150 2.6800 0.9600 2.1600 0.9600 2.1600 1.7800 1.7800 1.7800
                 1.7800 2.2000 1.6600 2.2000 1.6600 1.6600 2.0400 1.6600 2.0400 0.9600 1.9850 0.9600
                 1.9850 0.7500 1.7650 0.7500 1.7650 0.5000 1.8850 0.5000 1.8850 0.6300 2.1050 0.6300
                 2.1050 0.8400 2.8000 0.8400 ;
        POLYGON  1.9200 1.5400 1.6250 1.5400 1.6250 0.9900 0.2400 0.9900 0.2400 1.5550 0.5250 1.5550
                 0.5250 1.9200 0.4050 1.9200 0.4050 1.6750 0.1200 1.6750 0.1200 0.7500 0.3450 0.7500
                 0.3450 0.5000 0.4650 0.5000 0.4650 0.8700 1.7450 0.8700 1.7450 0.8800 1.8650 0.8800
                 1.8650 1.0000 1.7450 1.0000 1.7450 1.4200 1.9200 1.4200 ;
    END
END MX2X8

MACRO MX2X6
    CLASS CORE ;
    FOREIGN MX2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4100 1.5550 1.1700 1.6750 ;
        RECT  1.0500 1.3500 1.1700 1.6750 ;
        RECT  0.4100 1.1950 0.5300 1.6750 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0450 0.8500 1.4350 ;
        RECT  0.7300 1.0350 0.8500 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8700 1.2150 2.2500 1.4350 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.8700 1.2150 1.9900 1.4550 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2100 1.4300 4.3300 2.2100 ;
        RECT  3.9900 0.8000 4.2900 0.9200 ;
        RECT  4.1700 0.4050 4.2900 0.9200 ;
        RECT  4.0300 1.4300 4.3300 1.5500 ;
        RECT  4.0300 1.1900 4.1500 1.5500 ;
        RECT  3.3300 1.0400 4.1100 1.3100 ;
        RECT  3.9900 0.8000 4.1100 1.3100 ;
        RECT  3.3700 1.0400 3.4900 2.2100 ;
        RECT  3.3300 0.4050 3.4500 1.3100 ;
        RECT  2.6700 1.1900 4.1500 1.3100 ;
        RECT  2.6700 1.1750 2.8300 1.4350 ;
        RECT  2.5300 1.3600 2.7900 1.4800 ;
        RECT  2.6700 0.6300 2.7900 1.4800 ;
        RECT  2.4300 0.6300 2.7900 0.7500 ;
        RECT  2.5300 1.3600 2.6500 2.2100 ;
        RECT  2.4300 0.4000 2.5500 0.7500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  3.7500 -0.1800 3.8700 0.9200 ;
        RECT  2.9100 -0.1800 3.0300 0.9200 ;
        RECT  2.0100 -0.1800 2.1300 0.7400 ;
        RECT  0.7300 -0.1800 0.8500 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  3.7900 1.4300 3.9100 2.7900 ;
        RECT  2.9500 1.4300 3.0700 2.7900 ;
        RECT  2.1100 1.5550 2.2300 2.7900 ;
        RECT  0.5700 1.7950 0.6900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4900 1.2400 2.3700 1.2400 2.3700 0.9900 1.7500 0.9900 1.7500 1.8400 1.4300 1.8400
                 1.4300 2.2100 1.3100 2.2100 1.3100 1.7200 1.6300 1.7200 1.6300 0.9900 1.4700 0.9900
                 1.4700 0.6750 1.3700 0.6750 1.3700 0.4350 1.4900 0.4350 1.4900 0.5550 1.5900 0.5550
                 1.5900 0.8700 2.4900 0.8700 ;
        POLYGON  1.5100 1.6000 1.3900 1.6000 1.3900 1.2300 1.2300 1.2300 1.2300 0.9150 0.2400 0.9150
                 0.2400 1.5550 0.2700 1.5550 0.2700 2.0350 0.1500 2.0350 0.1500 1.6750 0.1200 1.6750
                 0.1200 0.6750 0.2500 0.6750 0.2500 0.5000 0.3700 0.5000 0.3700 0.7950 1.3500 0.7950
                 1.3500 1.1100 1.5100 1.1100 ;
    END
END MX2X6

MACRO MX2X4
    CLASS CORE ;
    FOREIGN MX2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.0600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9200 1.2000 1.2000 1.3200 ;
        RECT  0.3600 1.6000 1.0400 1.7200 ;
        RECT  0.9200 1.2000 1.0400 1.7200 ;
        RECT  0.3600 1.1750 0.5100 1.7200 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0250 0.8000 1.4800 ;
        RECT  0.6800 1.0000 0.8000 1.4800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.2300 2.3300 1.3950 ;
        RECT  1.8600 1.2750 2.1900 1.4050 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2400 1.4400 3.3600 2.2100 ;
        RECT  3.2200 0.5900 3.3400 0.8300 ;
        RECT  3.0600 1.4400 3.3600 1.5600 ;
        RECT  3.0400 0.7100 3.3400 0.8300 ;
        RECT  2.5600 1.3200 3.1800 1.4400 ;
        RECT  2.5600 0.7600 3.1600 0.8800 ;
        RECT  2.5600 1.1750 2.8300 1.4400 ;
        RECT  2.4000 1.5150 2.6800 1.6350 ;
        RECT  2.5600 0.6500 2.6800 1.6350 ;
        RECT  2.3200 0.6500 2.6800 0.7700 ;
        RECT  2.4000 1.5150 2.5200 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.0600 0.1800 ;
        RECT  3.6400 -0.1800 3.7600 0.6400 ;
        RECT  2.8000 -0.1800 2.9200 0.6400 ;
        RECT  1.9000 0.4600 2.1400 0.5800 ;
        RECT  1.9000 -0.1800 2.0200 0.5800 ;
        RECT  0.6800 -0.1800 0.8000 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.0600 2.7900 ;
        RECT  3.6600 1.5600 3.7800 2.7900 ;
        RECT  2.8200 1.5600 2.9400 2.7900 ;
        RECT  1.9800 1.5600 2.1000 2.7900 ;
        RECT  0.6400 1.8400 0.7600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4400 1.1100 1.7400 1.1100 1.7400 1.8400 1.4000 1.8400 1.4000 2.2100 1.2800 2.2100
                 1.2800 1.7200 1.6200 1.7200 1.6200 1.1100 1.5600 1.1100 1.5600 0.6400 1.3200 0.6400
                 1.3200 0.4000 1.4400 0.4000 1.4400 0.5200 1.6800 0.5200 1.6800 0.9900 2.4400 0.9900 ;
        POLYGON  1.5000 1.6000 1.3800 1.6000 1.3800 1.3500 1.3200 1.3500 1.3200 1.0000 1.1200 1.0000
                 1.1200 0.8800 0.2400 0.8800 0.2400 1.8400 0.3200 1.8400 0.3200 2.0800 0.2000 2.0800
                 0.2000 1.9600 0.1200 1.9600 0.1200 0.6400 0.2000 0.6400 0.2000 0.5000 0.3200 0.5000
                 0.3200 0.7600 1.4400 0.7600 1.4400 1.2300 1.5000 1.2300 ;
    END
END MX2X4

MACRO MX2X2
    CLASS CORE ;
    FOREIGN MX2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.6050 1.1850 1.7250 ;
        RECT  1.0650 1.3100 1.1850 1.7250 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6450 1.2800 0.8850 1.4850 ;
        RECT  0.6500 1.0900 0.8000 1.4850 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9050 1.2400 2.3050 1.3800 ;
        RECT  2.0450 1.2300 2.3050 1.3800 ;
        RECT  1.9050 1.2400 2.0250 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.1750 2.8300 1.4350 ;
        RECT  2.4250 1.1750 2.8300 1.2950 ;
        RECT  2.4250 0.5900 2.5450 1.6200 ;
        RECT  2.4050 1.5000 2.5250 2.2100 ;
        RECT  2.3450 0.4700 2.4650 0.7100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.7650 -0.1800 2.8850 0.6500 ;
        RECT  1.9250 -0.1800 2.0450 0.7100 ;
        RECT  0.6250 -0.1800 0.7450 0.7100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.8250 1.5600 2.9450 2.7900 ;
        RECT  1.9850 1.8500 2.1050 2.7900 ;
        RECT  0.7050 1.9700 0.8250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3050 1.1000 2.0650 1.1000 2.0650 0.9500 1.7850 0.9500 1.7850 2.0100 1.5250 2.0100
                 1.5250 2.0300 1.2850 2.0300 1.2850 1.9100 1.4050 1.9100 1.4050 1.8900 1.6650 1.8900
                 1.6650 0.9500 1.4250 0.9500 1.4250 0.7300 1.2650 0.7300 1.2650 0.4700 1.3850 0.4700
                 1.3850 0.6100 1.5450 0.6100 1.5450 0.8300 2.3050 0.8300 ;
        POLYGON  1.5450 1.7700 1.4250 1.7700 1.4250 1.1900 1.0650 1.1900 1.0650 0.9700 0.2400 0.9700
                 0.2400 1.8450 0.4050 1.8450 0.4050 2.0900 0.2850 2.0900 0.2850 1.9650 0.1200 1.9650
                 0.1200 0.7300 0.2050 0.7300 0.2050 0.4700 0.3250 0.4700 0.3250 0.8500 1.3050 0.8500
                 1.3050 1.0700 1.5450 1.0700 ;
    END
END MX2X2

MACRO MX2X1
    CLASS CORE ;
    FOREIGN MX2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.5800 1.1550 1.7000 ;
        RECT  1.0350 1.1200 1.1550 1.7000 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        RECT  0.3750 1.4600 0.4950 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0200 0.8150 1.4600 ;
        RECT  0.6950 1.0000 0.8150 1.4600 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.2100 2.0150 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3150 1.1750 2.5400 1.4350 ;
        RECT  2.3150 1.0550 2.4350 2.2100 ;
        RECT  2.2550 0.5900 2.3750 1.1750 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8350 -0.1800 1.9550 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8950 1.6000 2.0150 2.7900 ;
        RECT  0.5550 1.9200 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.1350 1.0900 1.6350 1.0900 1.6350 1.9400 1.3750 1.9400 1.3750 1.9800 1.1350 1.9800
                 1.1350 1.8600 1.2550 1.8600 1.2550 1.8200 1.5150 1.8200 1.5150 0.6400 1.1950 0.6400
                 1.1950 0.4000 1.3150 0.4000 1.3150 0.5200 1.6350 0.5200 1.6350 0.9700 2.1350 0.9700 ;
        POLYGON  1.3950 1.7000 1.2750 1.7000 1.2750 1.0000 1.0350 1.0000 1.0350 0.8800 0.2400 0.8800
                 0.2400 1.8450 0.2550 1.8450 0.2550 2.0850 0.1350 2.0850 0.1350 1.9650 0.1200 1.9650
                 0.1200 0.5200 0.1350 0.5200 0.1350 0.4000 0.2550 0.4000 0.2550 0.6400 0.2400 0.6400
                 0.2400 0.7600 1.3950 0.7600 ;
    END
END MX2X1

MACRO MDFFHQX8
    CLASS CORE ;
    FOREIGN MDFFHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 1.3450 2.7750 2.1900 ;
        RECT  2.6550 0.6650 2.7750 0.9850 ;
        RECT  2.6350 0.8650 2.7550 1.4650 ;
        RECT  0.0700 1.0250 2.7550 1.1450 ;
        RECT  1.8150 0.6650 1.9350 2.1900 ;
        RECT  0.9750 0.6650 1.0950 2.1850 ;
        RECT  0.1350 0.6650 0.2550 2.1850 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9450 1.1550 5.2050 1.3800 ;
        RECT  5.0850 0.9800 5.2050 1.3800 ;
        END
    END CK
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5350 1.2000 9.6550 1.4400 ;
        RECT  9.3500 1.2000 9.6550 1.4350 ;
        RECT  9.3500 1.1750 9.5000 1.4350 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7450 1.2100 11.1150 1.3950 ;
        RECT  10.7450 1.2100 11.0050 1.4200 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.2750 0.9700 11.3950 1.2100 ;
        RECT  11.0350 0.9400 11.2950 1.0900 ;
        RECT  10.2750 0.9700 11.3950 1.0900 ;
        RECT  10.0150 1.0000 10.3950 1.1200 ;
        RECT  10.0150 1.0000 10.1350 1.4400 ;
        END
    END S0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  11.0750 -0.1800 11.1950 0.8200 ;
        RECT  9.7950 -0.1800 9.9150 0.6400 ;
        RECT  7.4250 -0.1800 7.6650 0.3700 ;
        RECT  5.3250 -0.1800 5.5650 0.3800 ;
        RECT  3.9150 -0.1800 4.0350 0.6500 ;
        RECT  3.0750 -0.1800 3.1950 0.6500 ;
        RECT  2.2350 -0.1800 2.3550 0.6550 ;
        RECT  1.3950 -0.1800 1.5150 0.6550 ;
        RECT  0.5550 -0.1800 0.6750 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  10.9150 1.7800 11.0350 2.7900 ;
        RECT  9.5350 1.8500 9.6550 2.7900 ;
        RECT  7.4250 2.0700 7.6650 2.1900 ;
        RECT  7.4250 2.0700 7.5450 2.7900 ;
        RECT  5.6450 2.1000 5.7650 2.7900 ;
        RECT  3.9750 1.5400 4.0950 2.7900 ;
        RECT  3.0750 1.4450 3.1950 2.7900 ;
        RECT  2.2350 1.4450 2.3550 2.7900 ;
        RECT  1.3950 1.4450 1.5150 2.7900 ;
        RECT  0.5550 1.4450 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6350 1.6800 11.5550 1.6800 11.5550 1.8000 11.4350 1.8000 11.4350 1.6600
                 10.4150 1.6600 10.4150 1.2400 10.5350 1.2400 10.5350 1.5400 11.5150 1.5400
                 11.5150 0.8500 11.4950 0.8500 11.4950 0.5800 11.6150 0.5800 11.6150 0.7300
                 11.6350 0.7300 ;
        POLYGON  10.5550 0.8500 10.1550 0.8500 10.1550 0.8800 9.8950 0.8800 9.8950 1.5600
                 10.2950 1.5600 10.2950 2.2100 10.1750 2.2100 10.1750 1.6800 8.9850 1.6800
                 8.9850 1.7600 8.7450 1.7600 8.7450 1.5300 8.8650 1.5300 8.8650 0.7200 8.7850 0.7200
                 8.7850 0.6000 9.0250 0.6000 9.0250 0.7200 8.9850 0.7200 8.9850 1.5600 9.7750 1.5600
                 9.7750 0.7600 10.0350 0.7600 10.0350 0.7300 10.4350 0.7300 10.4350 0.5900
                 10.5550 0.5900 ;
        POLYGON  9.4350 0.8300 9.3150 0.8300 9.3150 0.4800 8.6650 0.4800 8.6650 1.1500 8.7050 1.1500
                 8.7050 1.3900 8.6650 1.3900 8.6650 1.4100 8.6250 1.4100 8.6250 1.8800 9.1750 1.8800
                 9.1750 2.0300 9.2950 2.0300 9.2950 2.1500 9.0550 2.1500 9.0550 2.0000 8.5050 2.0000
                 8.5050 1.2900 8.5450 1.2900 8.5450 0.4800 8.0650 0.4800 8.0650 0.8800 8.1450 0.8800
                 8.1450 1.1200 7.9450 1.1200 7.9450 0.6100 7.1850 0.6100 7.1850 0.4800 6.7050 0.4800
                 6.7050 0.9700 6.9650 0.9700 6.9650 1.2100 6.8450 1.2100 6.8450 1.0900 6.5850 1.0900
                 6.5850 0.3600 7.3050 0.3600 7.3050 0.4900 7.9450 0.4900 7.9450 0.3600 9.4350 0.3600 ;
        POLYGON  8.4250 0.7200 8.3850 0.7200 8.3850 1.9900 8.2650 1.9900 8.2650 1.3600 7.4650 1.3600
                 7.4650 1.3100 7.3250 1.3100 7.3250 1.1900 7.5850 1.1900 7.5850 1.2400 8.2650 1.2400
                 8.2650 0.7200 8.1850 0.7200 8.1850 0.6000 8.4250 0.6000 ;
        POLYGON  8.2250 2.2500 7.9850 2.2500 7.9850 1.9500 7.0450 1.9500 7.0450 2.2300 5.9250 2.2300
                 5.9250 0.8600 4.8250 0.8600 4.8250 1.5000 5.2450 1.5000 5.2450 1.7400 5.1250 1.7400
                 5.1250 1.6200 4.7050 1.6200 4.7050 0.6000 4.9650 0.6000 4.9650 0.7400 6.0450 0.7400
                 6.0450 2.1100 6.5850 2.1100 6.5850 1.3300 6.4250 1.3300 6.4250 1.2100 6.7050 1.2100
                 6.7050 2.1100 6.9250 2.1100 6.9250 1.8300 8.1050 1.8300 8.1050 2.1300 8.2250 2.1300 ;
        POLYGON  7.8250 1.1200 7.7050 1.1200 7.7050 1.0700 7.2050 1.0700 7.2050 1.4500 7.1250 1.4500
                 7.1250 1.7100 7.0050 1.7100 7.0050 1.3300 7.0850 1.3300 7.0850 0.8500 6.8250 0.8500
                 6.8250 0.6000 7.0650 0.6000 7.0650 0.7300 7.2050 0.7300 7.2050 0.9500 7.7050 0.9500
                 7.7050 0.8800 7.8250 0.8800 ;
        POLYGON  6.4650 1.9900 6.3450 1.9900 6.3450 1.5700 6.1850 1.5700 6.1850 0.6200 5.0850 0.6200
                 5.0850 0.4800 4.2750 0.4800 4.2750 1.1800 4.1550 1.1800 4.1550 0.3600 5.2050 0.3600
                 5.2050 0.5000 6.3050 0.5000 6.3050 1.4500 6.4650 1.4500 ;
        POLYGON  5.7250 1.9800 4.5150 1.9800 4.5150 2.1900 4.3950 2.1900 4.3950 1.4200 3.6750 1.4200
                 3.6750 2.1900 3.5550 2.1900 3.5550 1.5400 3.4950 1.5400 3.4950 1.2250 2.8750 1.2250
                 2.8750 1.1050 3.4950 1.1050 3.4950 0.6000 3.6150 0.6000 3.6150 1.3000 4.3950 1.3000
                 4.3950 0.6000 4.5150 0.6000 4.5150 1.8600 5.6050 1.8600 5.6050 1.1300 5.7250 1.1300 ;
    END
END MDFFHQX8

MACRO MDFFHQX4
    CLASS CORE ;
    FOREIGN MDFFHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1850 0.6300 2.3050 0.8700 ;
        RECT  1.9650 1.3150 2.2050 1.6500 ;
        RECT  2.0850 0.7500 2.2050 1.6500 ;
        RECT  1.2300 1.3150 2.2050 1.4350 ;
        RECT  1.3450 0.6300 1.4650 0.8700 ;
        RECT  1.0050 1.5300 1.3800 1.6500 ;
        RECT  1.2300 1.1750 1.3800 1.6500 ;
        RECT  1.2600 0.7500 1.3800 1.6500 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1750 0.6850 1.2950 ;
        RECT  0.5650 1.0550 0.6850 1.2950 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END CK
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5950 1.2000 7.7150 1.4400 ;
        RECT  7.3200 1.3150 7.7150 1.4350 ;
        RECT  7.3200 1.1750 7.4700 1.4350 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7150 1.2300 9.0600 1.4350 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0050 0.9900 9.3750 1.1100 ;
        RECT  8.2350 0.9700 9.2650 1.0900 ;
        RECT  9.0050 0.9400 9.2650 1.1100 ;
        RECT  8.0750 1.1900 8.3550 1.3100 ;
        RECT  8.2350 0.9700 8.3550 1.3100 ;
        RECT  8.0750 1.1900 8.1950 1.4400 ;
        END
    END S0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.1350 -0.1800 9.2550 0.8200 ;
        RECT  7.7550 -0.1800 7.8750 0.8300 ;
        RECT  5.4650 0.3900 5.7050 0.5100 ;
        RECT  5.5850 -0.1800 5.7050 0.5100 ;
        RECT  3.4450 -0.1800 3.5650 0.6800 ;
        RECT  2.6050 -0.1800 2.7250 0.6800 ;
        RECT  1.7650 -0.1800 1.8850 0.6800 ;
        RECT  0.9250 -0.1800 1.0450 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  8.9750 1.7950 9.0950 2.7900 ;
        RECT  7.5950 1.8500 7.7150 2.7900 ;
        RECT  5.4650 2.0700 5.7050 2.1900 ;
        RECT  5.4650 2.0700 5.5850 2.7900 ;
        RECT  3.4050 2.0100 3.6450 2.1300 ;
        RECT  3.4050 2.0100 3.5250 2.7900 ;
        RECT  2.4450 2.0100 2.6850 2.1300 ;
        RECT  2.4450 2.0100 2.5650 2.7900 ;
        RECT  1.4850 2.0100 1.7250 2.1300 ;
        RECT  1.4850 2.0100 1.6050 2.7900 ;
        RECT  0.5850 2.1100 0.7050 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.6750 0.8200 9.6150 0.8200 9.6150 1.6800 9.5750 1.6800 9.5750 1.8000 9.4550 1.8000
                 9.4550 1.6750 8.4750 1.6750 8.4750 1.2400 8.5950 1.2400 8.5950 1.5550 9.4950 1.5550
                 9.4950 0.7000 9.5550 0.7000 9.5550 0.5800 9.6750 0.5800 ;
        POLYGON  8.6150 0.8500 8.1150 0.8500 8.1150 1.0700 7.9550 1.0700 7.9550 1.5600 8.3550 1.5600
                 8.3550 2.2100 8.2350 2.2100 8.2350 1.6800 7.0250 1.6800 7.0250 1.7600 6.7850 1.7600
                 6.7850 1.5300 6.9050 1.5300 6.9050 0.7200 6.8850 0.7200 6.8850 0.6000 7.1250 0.6000
                 7.1250 0.7200 7.0250 0.7200 7.0250 1.5600 7.8350 1.5600 7.8350 0.9500 7.9950 0.9500
                 7.9950 0.7300 8.4950 0.7300 8.4950 0.5900 8.6150 0.5900 ;
        POLYGON  7.4550 0.8300 7.3350 0.8300 7.3350 0.4800 6.7650 0.4800 6.7650 1.3900 6.6650 1.3900
                 6.6650 1.8800 7.2350 1.8800 7.2350 2.0300 7.3550 2.0300 7.3550 2.1500 7.1150 2.1500
                 7.1150 2.0000 6.5450 2.0000 6.5450 1.1500 6.6450 1.1500 6.6450 0.4800 6.1650 0.4800
                 6.1650 0.8800 6.1850 0.8800 6.1850 1.1200 6.0450 1.1200 6.0450 0.7500 5.2250 0.7500
                 5.2250 0.4800 4.7450 0.4800 4.7450 1.0000 4.6650 1.0000 4.6650 1.2500 4.1250 1.2500
                 4.1250 1.3700 4.0050 1.3700 4.0050 1.1300 4.5450 1.1300 4.5450 0.8800 4.6250 0.8800
                 4.6250 0.3600 5.3450 0.3600 5.3450 0.6300 6.0450 0.6300 6.0450 0.3600 7.4550 0.3600 ;
        POLYGON  6.5250 0.7200 6.4250 0.7200 6.4250 1.9900 6.3050 1.9900 6.3050 1.3600 5.4850 1.3600
                 5.4850 1.3100 5.3650 1.3100 5.3650 1.1900 5.6050 1.1900 5.6050 1.2400 6.3050 1.2400
                 6.3050 0.7200 6.2850 0.7200 6.2850 0.6000 6.5250 0.6000 ;
        POLYGON  6.2650 2.2500 6.0250 2.2500 6.0250 1.9500 4.9250 1.9500 4.9250 2.2300 3.8450 2.2300
                 3.8450 1.8900 0.1350 1.8900 0.1350 1.6750 0.1200 1.6750 0.1200 0.9350 0.3250 0.9350
                 0.3250 0.6300 0.4450 0.6300 0.4450 1.0550 0.2400 1.0550 0.2400 1.5550 0.2550 1.5550
                 0.2550 1.7700 3.9650 1.7700 3.9650 2.1100 4.8050 2.1100 4.8050 1.2300 4.8850 1.2300
                 4.8850 1.1100 5.0050 1.1100 5.0050 1.3500 4.9250 1.3500 4.9250 1.8300 6.1450 1.8300
                 6.1450 2.1300 6.2650 2.1300 ;
        POLYGON  5.9250 1.0700 5.2450 1.0700 5.2450 1.5900 5.1650 1.5900 5.1650 1.7100 5.0450 1.7100
                 5.0450 1.4700 5.1250 1.4700 5.1250 0.9900 4.8650 0.9900 4.8650 0.6000 5.1050 0.6000
                 5.1050 0.8700 5.2450 0.8700 5.2450 0.9500 5.9250 0.9500 ;
        POLYGON  4.5050 0.7200 3.8850 0.7200 3.8850 1.4900 4.2450 1.4900 4.2450 1.4700 4.3650 1.4700
                 4.3650 1.9900 4.2450 1.9900 4.2450 1.6100 3.7650 1.6100 3.7650 1.3700 3.1850 1.3700
                 3.1850 1.1300 3.3050 1.1300 3.3050 1.2500 3.7650 1.2500 3.7650 0.6000 4.5050 0.6000 ;
        POLYGON  3.6450 1.1300 3.5250 1.1300 3.5250 1.0100 3.0650 1.0100 3.0650 1.5300 3.1650 1.5300
                 3.1650 1.6500 2.9250 1.6500 2.9250 1.5300 2.9450 1.5300 2.9450 1.0100 2.5450 1.0100
                 2.5450 1.1900 2.4250 1.1900 2.4250 0.8900 2.9450 0.8900 2.9450 0.6600 3.0250 0.6600
                 3.0250 0.5400 3.1450 0.5400 3.1450 0.8900 3.6450 0.8900 ;
    END
END MDFFHQX4

MACRO MDFFHQX2
    CLASS CORE ;
    FOREIGN MDFFHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.4650 1.3350 1.5850 ;
        RECT  1.2150 1.3450 1.3350 1.5850 ;
        RECT  0.9400 1.4650 1.0900 1.7250 ;
        END
    END CK
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4850 0.9600 6.6800 1.2000 ;
        RECT  6.4500 0.8850 6.6750 1.1450 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9000 1.0250 8.0600 1.4800 ;
        RECT  7.9400 1.0000 8.0600 1.4800 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4250 1.2300 8.6850 1.3800 ;
        RECT  8.4250 1.0700 8.5450 1.3800 ;
        RECT  8.3400 0.7600 8.4600 1.1900 ;
        RECT  8.2200 1.0700 8.5450 1.1900 ;
        RECT  7.3000 0.7600 8.4600 0.8800 ;
        RECT  7.5400 0.7600 7.7800 1.0900 ;
        RECT  7.0400 1.0000 7.4200 1.1200 ;
        RECT  7.3000 0.7600 7.4200 1.1200 ;
        RECT  7.0400 1.0000 7.1600 1.4400 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6800 0.6750 2.2050 ;
        RECT  0.3600 1.1750 0.6750 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.1000 -0.1800 8.2200 0.6400 ;
        RECT  6.8200 -0.1800 6.9400 0.6400 ;
        RECT  4.4300 0.3800 4.6700 0.5000 ;
        RECT  4.5500 -0.1800 4.6700 0.5000 ;
        RECT  2.5700 -0.1800 2.6900 0.6800 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  7.9400 1.8400 8.0600 2.7900 ;
        RECT  6.5600 1.5600 6.6800 2.7900 ;
        RECT  4.4300 2.0600 4.6700 2.1800 ;
        RECT  4.4300 2.0600 4.5500 2.7900 ;
        RECT  2.3100 2.0600 2.4300 2.7900 ;
        RECT  0.9750 1.8450 1.0950 2.7900 ;
        RECT  0.1350 1.5550 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.9250 1.7200 8.5400 1.7200 8.5400 1.8400 8.4200 1.8400 8.4200 1.7200 7.4400 1.7200
                 7.4400 1.2400 7.5600 1.2400 7.5600 1.6000 8.8050 1.6000 8.8050 0.9500 8.5800 0.9500
                 8.5800 0.5900 8.7000 0.5900 8.7000 0.8300 8.9250 0.8300 ;
        POLYGON  7.5800 0.6400 7.1800 0.6400 7.1800 0.8800 6.9200 0.8800 6.9200 1.5600 7.3200 1.5600
                 7.3200 2.2100 7.2000 2.2100 7.2000 1.6800 6.8000 1.6800 6.8000 1.4400 5.9900 1.4400
                 5.9900 1.5800 5.9500 1.5800 5.9500 1.7000 5.8300 1.7000 5.8300 1.4600 5.8700 1.4600
                 5.8700 0.7200 5.8300 0.7200 5.8300 0.6000 6.0700 0.6000 6.0700 0.7200 5.9900 0.7200
                 5.9900 1.3200 6.8000 1.3200 6.8000 0.7600 7.0600 0.7600 7.0600 0.5200 7.4600 0.5200
                 7.4600 0.4000 7.5800 0.4000 ;
        POLYGON  6.4600 0.6600 6.3400 0.6600 6.3400 0.4800 5.7100 0.4800 5.7100 1.1000 5.7500 1.1000
                 5.7500 1.3400 5.7100 1.3400 5.7100 1.9100 6.2600 1.9100 6.2600 2.0300 5.5900 2.0300
                 5.5900 0.4800 5.1100 0.4800 5.1100 0.9200 5.2300 0.9200 5.2300 1.0400 4.9900 1.0400
                 4.9900 0.7400 4.1900 0.7400 4.1900 0.4800 3.7100 0.4800 3.7100 0.9800 3.5700 0.9800
                 3.5700 1.2600 2.9900 1.2600 2.9900 1.3800 2.8700 1.3800 2.8700 1.1400 3.4500 1.1400
                 3.4500 0.8600 3.5900 0.8600 3.5900 0.3600 4.3100 0.3600 4.3100 0.6200 4.9900 0.6200
                 4.9900 0.3600 6.4600 0.3600 ;
        POLYGON  5.4700 1.9800 5.3500 1.9800 5.3500 1.3000 4.2900 1.3000 4.2900 1.1800 5.3500 1.1800
                 5.3500 0.7200 5.2300 0.7200 5.2300 0.6000 5.4700 0.6000 ;
        POLYGON  5.2500 2.2400 5.0100 2.2400 5.0100 1.9400 3.8900 1.9400 3.8900 2.2200 2.7100 2.2200
                 2.7100 1.9400 2.0350 1.9400 2.0350 1.9650 1.5150 1.9650 1.5150 2.0850 1.3950 2.0850
                 1.3950 1.8450 1.4550 1.8450 1.4550 0.6800 1.5750 0.6800 1.5750 1.8450 1.9150 1.8450
                 1.9150 1.8200 2.8300 1.8200 2.8300 2.1000 3.7700 2.1000 3.7700 1.2200 3.8100 1.2200
                 3.8100 1.1000 3.9300 1.1000 3.9300 1.3400 3.8900 1.3400 3.8900 1.8200 5.1300 1.8200
                 5.1300 2.1200 5.2500 2.1200 ;
        POLYGON  4.8700 1.0600 4.1700 1.0600 4.1700 1.5800 4.1300 1.5800 4.1300 1.7000 4.0100 1.7000
                 4.0100 1.4600 4.0500 1.4600 4.0500 0.9800 3.8300 0.9800 3.8300 0.6000 4.0700 0.6000
                 4.0700 0.8600 4.1700 0.8600 4.1700 0.9400 4.8700 0.9400 ;
        POLYGON  3.4700 0.7200 2.9300 0.7200 2.9300 1.0200 2.7500 1.0200 2.7500 1.5000 3.1100 1.5000
                 3.1100 1.4600 3.2300 1.4600 3.2300 1.9800 3.1100 1.9800 3.1100 1.6200 2.0700 1.6200
                 2.0700 1.3400 2.0500 1.3400 2.0500 1.1000 2.1900 1.1000 2.1900 1.5000 2.6300 1.5000
                 2.6300 0.9000 2.8100 0.9000 2.8100 0.6000 3.4700 0.6000 ;
        POLYGON  2.5100 1.3800 2.3900 1.3800 2.3900 0.9800 1.9300 0.9800 1.9300 1.4600 1.9500 1.4600
                 1.9500 1.7000 1.8300 1.7000 1.8300 1.5800 1.8100 1.5800 1.8100 0.5600 1.3350 0.5600
                 1.3350 1.1800 0.7950 1.1800 0.7950 1.0600 1.2150 1.0600 1.2150 0.4400 2.2700 0.4400
                 2.2700 0.8600 2.5100 0.8600 ;
    END
END MDFFHQX2

MACRO MDFFHQX1
    CLASS CORE ;
    FOREIGN MDFFHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7100 1.0900 0.8600 1.4250 ;
        RECT  0.6500 1.0950 0.8300 1.4350 ;
        END
    END CK
    PIN D0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0650 0.9600 6.1850 1.2000 ;
        RECT  5.8700 0.9600 6.1850 1.1450 ;
        RECT  5.8700 0.8850 6.0200 1.1450 ;
        END
    END D0
    PIN D1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.2100 7.6250 1.4100 ;
        RECT  7.2650 1.2100 7.5250 1.4350 ;
        END
    END D1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7650 0.9700 7.8850 1.2100 ;
        RECT  7.5550 0.9400 7.8150 1.0900 ;
        RECT  6.5450 0.9700 7.8850 1.0900 ;
        RECT  6.5450 0.9700 6.6650 1.4400 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.2950 0.2650 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.6650 -0.1800 7.7850 0.8200 ;
        RECT  6.0650 -0.1800 6.1850 0.6400 ;
        RECT  3.7950 0.3900 4.0350 0.5100 ;
        RECT  3.7950 -0.1800 3.9150 0.5100 ;
        RECT  2.0150 -0.1800 2.1350 0.6800 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.4450 1.7950 7.5650 2.7900 ;
        RECT  6.0650 1.5600 6.1850 2.7900 ;
        RECT  3.7950 2.0700 4.0350 2.1900 ;
        RECT  3.7950 2.0700 3.9150 2.7900 ;
        RECT  1.7150 2.0100 1.9550 2.1300 ;
        RECT  1.7150 2.0100 1.8350 2.7900 ;
        RECT  0.5650 1.8500 0.6850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.2050 0.8200 8.1250 0.8200 8.1250 1.6800 8.0450 1.6800 8.0450 1.8000 7.9250 1.8000
                 7.9250 1.6750 6.9450 1.6750 6.9450 1.2400 7.0650 1.2400 7.0650 1.5550 8.0050 1.5550
                 8.0050 0.7000 8.0850 0.7000 8.0850 0.5800 8.2050 0.5800 ;
        POLYGON  7.1450 0.8500 6.4250 0.8500 6.4250 1.5600 6.8250 1.5600 6.8250 2.2100 6.7050 2.2100
                 6.7050 1.6800 6.3050 1.6800 6.3050 1.4400 5.3550 1.4400 5.3550 1.5900 5.2550 1.5900
                 5.2550 1.9900 5.1350 1.9900 5.1350 1.4700 5.2350 1.4700 5.2350 0.7200 5.1350 0.7200
                 5.1350 0.6000 5.3750 0.6000 5.3750 0.7200 5.3550 0.7200 5.3550 1.3200 6.3050 1.3200
                 6.3050 0.7300 7.0250 0.7300 7.0250 0.5900 7.1450 0.5900 ;
        POLYGON  5.7650 1.8600 5.6450 1.8600 5.6450 1.9800 5.4950 1.9800 5.4950 2.2300 4.8950 2.2300
                 4.8950 0.4800 4.4150 0.4800 4.4150 0.8400 4.5350 0.8400 4.5350 1.1000 4.4150 1.1000
                 4.4150 0.9600 4.2950 0.9600 4.2950 0.7500 3.5550 0.7500 3.5550 0.4800 3.0750 0.4800
                 3.0750 0.9800 3.0350 0.9800 3.0350 1.1000 3.0150 1.1000 3.0150 1.2700 2.4550 1.2700
                 2.4550 1.3900 2.3350 1.3900 2.3350 1.1500 2.8950 1.1500 2.8950 0.8600 2.9550 0.8600
                 2.9550 0.3600 3.6750 0.3600 3.6750 0.6300 4.2950 0.6300 4.2950 0.3600 5.7050 0.3600
                 5.7050 0.8100 5.5850 0.8100 5.5850 0.4800 5.0150 0.4800 5.0150 1.1100 5.1150 1.1100
                 5.1150 1.3500 5.0150 1.3500 5.0150 2.1100 5.3750 2.1100 5.3750 1.8600 5.5250 1.8600
                 5.5250 1.7400 5.7650 1.7400 ;
        POLYGON  4.7750 1.9900 4.6550 1.9900 4.6550 1.5600 3.7550 1.5600 3.7550 1.1300 3.8750 1.1300
                 3.8750 1.4400 4.6550 1.4400 4.6550 0.7200 4.5350 0.7200 4.5350 0.6000 4.7750 0.6000 ;
        POLYGON  4.5950 2.2500 4.3550 2.2500 4.3550 1.9500 3.2550 1.9500 3.2550 2.2300 2.0750 2.2300
                 2.0750 1.8900 1.1050 1.8900 1.1050 2.1000 0.9850 2.1000 0.9850 1.2900 1.0350 1.2900
                 1.0350 0.6800 1.1550 0.6800 1.1550 1.4100 1.1050 1.4100 1.1050 1.7700 2.1950 1.7700
                 2.1950 2.1100 3.1350 2.1100 3.1350 1.2300 3.2750 1.2300 3.2750 1.1100 3.3950 1.1100
                 3.3950 1.3500 3.2550 1.3500 3.2550 1.8300 4.4750 1.8300 4.4750 2.1300 4.5950 2.1300 ;
        POLYGON  4.1950 1.3200 4.0550 1.3200 4.0550 1.0100 3.6350 1.0100 3.6350 1.5900 3.4950 1.5900
                 3.4950 1.7100 3.3750 1.7100 3.3750 1.4700 3.5150 1.4700 3.5150 0.9900 3.1950 0.9900
                 3.1950 0.6000 3.4350 0.6000 3.4350 0.8700 3.6350 0.8700 3.6350 0.8900 4.1750 0.8900
                 4.1750 1.0800 4.1950 1.0800 ;
        POLYGON  2.8350 0.7200 2.3750 0.7200 2.3750 1.0300 2.2150 1.0300 2.2150 1.5100 2.5750 1.5100
                 2.5750 1.4700 2.6950 1.4700 2.6950 1.9900 2.5750 1.9900 2.5750 1.6300 1.5950 1.6300
                 1.5950 1.3700 1.5150 1.3700 1.5150 1.1300 1.7150 1.1300 1.7150 1.5100 2.0950 1.5100
                 2.0950 0.9100 2.2550 0.9100 2.2550 0.6000 2.8350 0.6000 ;
        POLYGON  1.9750 1.3900 1.8550 1.3900 1.8550 1.0100 1.3950 1.0100 1.3950 1.5300 1.4750 1.5300
                 1.4750 1.6500 1.2350 1.6500 1.2350 1.5300 1.2750 1.5300 1.2750 0.5600 0.9150 0.5600
                 0.9150 0.9700 0.5200 0.9700 0.5200 1.2400 0.4000 1.2400 0.4000 0.8500 0.7950 0.8500
                 0.7950 0.4400 1.7150 0.4400 1.7150 0.8900 1.9750 0.8900 ;
    END
END MDFFHQX1

MACRO INVXL
    CLASS CORE ;
    FOREIGN INVXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.8700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 1.0400 0.2400 1.4550 ;
        RECT  0.0700 1.0400 0.2400 1.4450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6800 0.6750 1.6950 ;
        RECT  0.3600 1.1750 0.6750 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.8700 0.1800 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.8700 2.7900 ;
        RECT  0.1350 1.5750 0.2550 2.7900 ;
        END
    END VDD
END INVXL

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9050 1.2050 2.2650 1.3250 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1450 0.7400 3.3850 0.8600 ;
        RECT  3.2050 1.4700 3.3250 2.2100 ;
        RECT  0.7450 0.7900 3.2650 0.9100 ;
        RECT  0.6850 1.5000 3.3250 1.6200 ;
        RECT  2.3850 0.7900 2.5400 1.1450 ;
        RECT  2.3850 0.7900 2.5050 1.6200 ;
        RECT  2.3650 1.4700 2.4850 2.2100 ;
        RECT  2.3650 0.6700 2.4850 0.9100 ;
        RECT  1.4650 0.7400 1.7050 0.9100 ;
        RECT  1.5250 1.4650 1.6450 2.2100 ;
        RECT  0.6250 0.7400 0.8650 0.8600 ;
        RECT  0.6850 1.5000 0.8050 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.7850 -0.1800 2.9050 0.6700 ;
        RECT  1.9450 -0.1800 2.0650 0.6700 ;
        RECT  1.1050 -0.1800 1.2250 0.6700 ;
        RECT  0.2650 -0.1800 0.3850 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.7850 1.7400 2.9050 2.7900 ;
        RECT  1.9450 1.7400 2.0650 2.7900 ;
        RECT  1.1050 1.7400 1.2250 2.7900 ;
        RECT  0.2650 1.4650 0.3850 2.7900 ;
        END
    END VDD
END INVX8

MACRO INVX6
    CLASS CORE ;
    FOREIGN INVX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8400 1.1500 1.4000 1.2700 ;
        RECT  0.8850 1.1500 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3200 1.4300 2.4400 2.2100 ;
        RECT  0.5800 0.9100 2.4400 1.0300 ;
        RECT  2.3200 0.4000 2.4400 1.0300 ;
        RECT  0.6400 1.5000 2.4400 1.6200 ;
        RECT  1.5200 1.1750 1.6700 1.6200 ;
        RECT  1.5200 0.9100 1.6400 1.6200 ;
        RECT  1.4800 1.4300 1.6000 2.2100 ;
        RECT  1.4800 0.4000 1.6000 1.0300 ;
        RECT  0.6400 1.4300 0.7600 2.2100 ;
        RECT  0.5800 0.4000 0.7000 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.9000 -0.1800 2.0200 0.7900 ;
        RECT  1.0600 -0.1800 1.1800 0.7900 ;
        RECT  0.1600 -0.1800 0.2800 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.9000 1.7400 2.0200 2.7900 ;
        RECT  1.0600 1.7400 1.1800 2.7900 ;
        RECT  0.2200 1.4300 0.3400 2.7900 ;
        END
    END VDD
END INVX6

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8000 1.2600 1.4000 1.3800 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.5200 0.8500 1.6400 1.7250 ;
        RECT  1.5000 1.5000 1.6200 2.2100 ;
        RECT  0.6600 0.8500 1.6400 0.9700 ;
        RECT  1.5000 0.6800 1.6200 0.9700 ;
        RECT  0.6600 1.5000 1.6700 1.6200 ;
        RECT  0.6600 1.5000 0.7800 2.2100 ;
        RECT  0.6600 0.6800 0.7800 0.9700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.9200 -0.1800 2.0400 0.7300 ;
        RECT  1.0800 -0.1800 1.2000 0.7300 ;
        RECT  0.2400 -0.1800 0.3600 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.9200 1.5600 2.0400 2.7900 ;
        RECT  1.0800 1.7400 1.2000 2.7900 ;
        RECT  0.2400 1.5600 0.3600 2.7900 ;
        END
    END VDD
END INVX4

MACRO INVX3
    CLASS CORE ;
    FOREIGN INVX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3240  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.7900 0.4150 1.2450 ;
        RECT  0.2950 0.7600 0.4150 1.2450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.1250 1.5150 2.0150 ;
        RECT  0.6500 0.7600 1.5150 0.8800 ;
        RECT  1.3950 0.5900 1.5150 0.8800 ;
        RECT  0.6500 1.1250 1.5150 1.2450 ;
        RECT  0.6500 0.7600 0.8000 1.2450 ;
        RECT  0.6500 0.7100 0.7700 1.4850 ;
        RECT  0.5550 1.3650 0.6750 2.0150 ;
        RECT  0.5550 0.5900 0.6750 0.8300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.3650 1.0950 2.7900 ;
        RECT  0.1350 1.3650 0.2550 2.7900 ;
        END
    END VDD
END INVX3

MACRO INVX20
    CLASS CORE ;
    FOREIGN INVX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.1600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 1.1650 6.3650 1.2850 ;
        RECT  0.8850 1.1650 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.6132  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2850 1.4500 7.4050 2.2100 ;
        RECT  0.5550 0.9250 7.4050 1.0450 ;
        RECT  7.2850 0.4000 7.4050 1.0450 ;
        RECT  0.5650 1.5000 7.4050 1.6200 ;
        RECT  6.7400 1.1750 6.8900 1.6200 ;
        RECT  6.4850 1.3150 6.8900 1.6200 ;
        RECT  6.4850 0.9250 6.6050 1.6200 ;
        RECT  6.4450 1.4450 6.5650 2.2100 ;
        RECT  6.4450 0.4000 6.5650 1.0450 ;
        RECT  5.6050 1.4450 5.7250 2.2100 ;
        RECT  5.6050 0.4000 5.7250 1.0450 ;
        RECT  4.7650 1.4450 4.8850 2.2100 ;
        RECT  4.7650 0.4000 4.8850 1.0450 ;
        RECT  3.9250 1.4450 4.0450 2.2100 ;
        RECT  3.9250 0.4000 4.0450 1.0450 ;
        RECT  3.0850 1.4450 3.2050 2.2100 ;
        RECT  3.0850 0.4000 3.2050 1.0450 ;
        RECT  2.2450 1.4450 2.3650 2.2100 ;
        RECT  2.2450 0.4000 2.3650 1.0450 ;
        RECT  1.4050 1.4450 1.5250 2.2100 ;
        RECT  1.3950 0.4000 1.5150 1.0450 ;
        RECT  0.5650 1.4450 0.6850 2.2100 ;
        RECT  0.5550 0.4000 0.6750 1.0450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.8650 -0.1800 6.9850 0.8050 ;
        RECT  6.0250 -0.1800 6.1450 0.8050 ;
        RECT  5.1850 -0.1800 5.3050 0.8050 ;
        RECT  4.3450 -0.1800 4.4650 0.8050 ;
        RECT  3.5050 -0.1800 3.6250 0.8050 ;
        RECT  2.6650 -0.1800 2.7850 0.8050 ;
        RECT  1.8250 -0.1800 1.9450 0.8050 ;
        RECT  0.9750 -0.1800 1.0950 0.8050 ;
        RECT  0.1350 -0.1800 0.2550 0.9100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.8650 1.7400 6.9850 2.7900 ;
        RECT  6.0250 1.7400 6.1450 2.7900 ;
        RECT  5.1850 1.7400 5.3050 2.7900 ;
        RECT  4.3450 1.7400 4.4650 2.7900 ;
        RECT  3.5050 1.7400 3.6250 2.7900 ;
        RECT  2.6650 1.7400 2.7850 2.7900 ;
        RECT  1.8250 1.7400 1.9450 2.7900 ;
        RECT  0.9850 1.7400 1.1050 2.7900 ;
        RECT  0.1450 1.4450 0.2650 2.7900 ;
        END
    END VDD
END INVX20

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.4500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3700 1.0000 0.4900 1.2400 ;
        RECT  0.0700 1.0250 0.4900 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        RECT  0.6500 0.6800 0.7700 2.0100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.4500 0.1800 ;
        RECT  1.0700 -0.1800 1.1900 0.7300 ;
        RECT  0.2300 -0.1800 0.3500 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.4500 2.7900 ;
        RECT  1.0700 1.3600 1.1900 2.7900 ;
        RECT  0.2300 1.3600 0.3500 2.7900 ;
        END
    END VDD
END INVX2

MACRO INVX16
    CLASS CORE ;
    FOREIGN INVX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.7280  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.2050 5.4950 1.3250 ;
        RECT  0.8850 1.2050 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5000 5.7350 1.6200 ;
        RECT  5.6150 0.7900 5.7350 1.6200 ;
        RECT  5.5800 1.4650 5.7300 1.7250 ;
        RECT  5.5950 1.4650 5.7150 2.2100 ;
        RECT  0.6150 0.7900 5.7350 0.9100 ;
        RECT  5.5950 0.6700 5.7150 0.9100 ;
        RECT  4.6950 0.7400 4.9350 0.9100 ;
        RECT  4.7550 1.4700 4.8750 2.2100 ;
        RECT  3.8550 0.7400 4.0950 0.9100 ;
        RECT  3.9150 1.4700 4.0350 2.2100 ;
        RECT  3.0150 0.7400 3.2550 0.9100 ;
        RECT  3.0750 1.4650 3.1950 2.2100 ;
        RECT  2.1750 0.7400 2.4150 0.9100 ;
        RECT  2.2350 1.4650 2.3550 2.2100 ;
        RECT  1.3350 0.7400 1.5750 0.9100 ;
        RECT  1.3950 1.4650 1.5150 2.2100 ;
        RECT  0.4950 0.7400 0.7350 0.8600 ;
        RECT  0.5550 1.4650 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  6.0150 -0.1800 6.1350 0.6700 ;
        RECT  5.1750 -0.1800 5.2950 0.6700 ;
        RECT  4.3350 -0.1800 4.4550 0.6700 ;
        RECT  3.4950 -0.1800 3.6150 0.6700 ;
        RECT  2.6550 -0.1800 2.7750 0.6700 ;
        RECT  1.8150 -0.1800 1.9350 0.6700 ;
        RECT  0.9750 -0.1800 1.0950 0.6650 ;
        RECT  0.1350 -0.1800 0.2550 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  6.0150 1.4700 6.1350 2.7900 ;
        RECT  5.1750 1.7400 5.2950 2.7900 ;
        RECT  4.3350 1.7400 4.4550 2.7900 ;
        RECT  3.4950 1.7400 3.6150 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.4650 0.2550 2.7900 ;
        END
    END VDD
END INVX16

MACRO INVX12
    CLASS CORE ;
    FOREIGN INVX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.2960  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 1.1500 3.8350 1.2700 ;
        RECT  0.8850 1.1500 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5000 4.0750 1.6200 ;
        RECT  3.9550 0.9100 4.0750 1.6200 ;
        RECT  3.9150 1.4300 4.0350 2.2100 ;
        RECT  0.5550 0.9100 4.0750 1.0300 ;
        RECT  3.9150 0.4000 4.0350 1.0300 ;
        RECT  3.8400 1.4650 4.0350 1.7250 ;
        RECT  3.0750 1.4300 3.1950 2.2100 ;
        RECT  3.0750 0.4000 3.1950 1.0300 ;
        RECT  2.2350 1.4300 2.3550 2.2100 ;
        RECT  2.2350 0.4000 2.3550 1.0300 ;
        RECT  1.3950 1.4300 1.5150 2.2100 ;
        RECT  1.3950 0.4000 1.5150 1.0300 ;
        RECT  0.5550 1.4300 0.6750 2.2100 ;
        RECT  0.5550 0.4000 0.6750 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  4.3350 -0.1800 4.4550 0.9150 ;
        RECT  3.4950 -0.1800 3.6150 0.7900 ;
        RECT  2.6550 -0.1800 2.7750 0.7900 ;
        RECT  1.8150 -0.1800 1.9350 0.7900 ;
        RECT  0.9750 -0.1800 1.0950 0.7900 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  4.3350 1.4300 4.4550 2.7900 ;
        RECT  3.4950 1.7400 3.6150 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.4300 0.2550 2.7900 ;
        END
    END VDD
END INVX12

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.8700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 0.7950 0.2400 1.2200 ;
        RECT  0.0700 0.7950 0.2400 1.2000 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6250 0.6750 1.9900 ;
        RECT  0.3600 0.8850 0.6750 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.8700 0.1800 ;
        RECT  0.1350 -0.1800 0.2550 0.6750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.8700 2.7900 ;
        RECT  0.1350 1.3400 0.2550 2.7900 ;
        END
    END VDD
END INVX1

MACRO HOLDX1
    CLASS CORE ;
    FOREIGN HOLDX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4850 0.6800 1.6050 1.6000 ;
        RECT  0.4050 1.3600 1.6050 1.4800 ;
        RECT  1.2300 1.1750 1.6050 1.4800 ;
        RECT  0.4050 1.0200 0.5250 1.4800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  0.8850 1.2400 0.7650 1.2400 0.7650 0.9000 0.2550 0.9000 0.2550 1.9900 0.1350 1.9900
                 0.1350 0.6600 0.2550 0.6600 0.2550 0.7800 0.8850 0.7800 ;
    END
END HOLDX1

MACRO FILL8
    CLASS CORE ;
    FOREIGN FILL8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        END
    END VSS
END FILL8

MACRO FILL64
    CLASS CORE ;
    FOREIGN FILL64 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 18.5600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 18.5600 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 18.5600 0.1800 ;
        END
    END VSS
END FILL64

MACRO FILL4
    CLASS CORE ;
    FOREIGN FILL4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.1600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.1600 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.1600 0.1800 ;
        END
    END VSS
END FILL4

MACRO FILL32
    CLASS CORE ;
    FOREIGN FILL32 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        END
    END VSS
END FILL32

MACRO FILL2
    CLASS CORE ;
    FOREIGN FILL2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.5800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.5800 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.5800 0.1800 ;
        END
    END VSS
END FILL2

MACRO FILL16
    CLASS CORE ;
    FOREIGN FILL16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        END
    END VSS
END FILL16

MACRO FILL1
    CLASS CORE ;
    FOREIGN FILL1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.2900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.2900 0.1800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.2900 2.7900 ;
        END
    END VDD
END FILL1

MACRO EDFFXL
    CLASS CORE ;
    FOREIGN EDFFXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1300 0.5100 1.6000 ;
        RECT  0.3800 1.1300 0.5000 1.6300 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3900 1.1950 6.6550 1.4450 ;
        RECT  6.3950 1.1750 6.6550 1.4450 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0300 1.1750 7.1800 1.4350 ;
        RECT  6.8900 1.1950 7.1800 1.4350 ;
        RECT  5.7700 1.5650 6.9700 1.6850 ;
        RECT  6.8500 1.3150 6.9700 1.6850 ;
        RECT  5.2700 2.1300 5.8900 2.2500 ;
        RECT  5.7700 0.9600 5.8900 2.2500 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5400 0.7400 7.7800 0.8600 ;
        RECT  7.6100 0.7400 7.7600 1.1450 ;
        RECT  7.6000 1.0050 7.7200 1.5800 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3150 0.6800 9.4350 2.0900 ;
        RECT  9.0600 1.4650 9.4350 1.7250 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.8950 -0.1800 9.0150 0.9200 ;
        RECT  8.0800 -0.1800 8.2000 0.4000 ;
        RECT  6.6100 0.4550 6.8500 0.5750 ;
        RECT  6.6100 -0.1800 6.7300 0.5750 ;
        RECT  4.5900 0.6800 4.8300 0.8000 ;
        RECT  4.5900 -0.1800 4.7100 0.8000 ;
        RECT  2.5700 0.6000 2.8100 0.7200 ;
        RECT  2.5700 -0.1800 2.6900 0.7200 ;
        RECT  0.5600 -0.1800 0.6800 0.7700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.8950 1.9700 9.0150 2.7900 ;
        RECT  8.0800 1.9800 8.2000 2.7900 ;
        RECT  6.6100 1.8050 6.8500 1.9250 ;
        RECT  6.6100 1.8050 6.7300 2.7900 ;
        RECT  4.5900 2.2300 4.7100 2.7900 ;
        RECT  2.6900 2.0400 2.8100 2.7900 ;
        RECT  2.5700 2.0400 2.8100 2.1600 ;
        RECT  0.5600 1.7500 0.6800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.1950 1.3400 8.6800 1.3400 8.6800 1.5800 8.5600 1.5800 8.5600 0.9200 8.5050 0.9200
                 8.5050 0.6800 8.6250 0.6800 8.6250 0.8000 8.6800 0.8000 8.6800 1.2200 9.1950 1.2200 ;
        POLYGON  7.9400 0.5200 7.4500 0.5200 7.4500 0.5000 7.0900 0.5000 7.0900 0.8150 6.1750 0.8150
                 6.1750 0.5000 5.1900 0.5000 5.1900 0.8600 5.1700 0.8600 5.1700 1.6500 5.2500 1.6500
                 5.2500 1.7700 5.0100 1.7700 5.0100 1.6500 5.0500 1.6500 5.0500 1.4900 4.4300 1.4900
                 4.4300 1.2500 4.5500 1.2500 4.5500 1.3700 5.0500 1.3700 5.0500 0.7400 5.0700 0.7400
                 5.0700 0.3800 6.2950 0.3800 6.2950 0.6950 6.9700 0.6950 6.9700 0.3800 7.5700 0.3800
                 7.5700 0.4000 7.9400 0.4000 ;
        POLYGON  7.4200 1.7700 7.0900 1.7700 7.0900 1.6500 7.3000 1.6500 7.3000 1.0550 6.2300 1.0550
                 6.2300 1.4400 6.1100 1.4400 6.1100 0.9350 7.2100 0.9350 7.2100 0.6200 7.3300 0.6200
                 7.3300 0.8150 7.4200 0.8150 ;
        POLYGON  5.6500 2.0100 4.3000 2.0100 4.3000 2.0900 3.6500 2.0900 3.6500 2.0100 3.1700 2.0100
                 3.1700 1.6800 2.2100 1.6800 2.2100 2.0100 1.4900 2.0100 1.4900 1.9500 1.3700 1.9500
                 1.3700 0.6200 1.4900 0.6200 1.4900 1.8300 1.6100 1.8300 1.6100 1.8900 2.0900 1.8900
                 2.0900 1.5600 3.2900 1.5600 3.2900 1.8900 3.7700 1.8900 3.7700 1.9700 4.1800 1.9700
                 4.1800 1.8900 5.5300 1.8900 5.5300 0.6200 5.6500 0.6200 ;
        POLYGON  4.9300 1.2500 4.8100 1.2500 4.8100 1.1300 4.3100 1.1300 4.3100 1.7300 4.0100 1.7300
                 4.0100 1.8500 3.8900 1.8500 3.8900 1.6100 4.1900 1.6100 4.1900 1.1300 3.8900 1.1300
                 3.8900 0.6200 4.0100 0.6200 4.0100 1.0100 4.9300 1.0100 ;
        POLYGON  4.0700 1.4900 3.9500 1.4900 3.9500 1.3700 3.6500 1.3700 3.6500 1.2000 3.4100 1.2000
                 3.4100 0.9600 3.6500 0.9600 3.6500 0.5600 3.0500 0.5600 3.0500 0.9600 2.3300 0.9600
                 2.3300 0.5000 1.7300 0.5000 1.7300 1.4900 1.6100 1.4900 1.6100 0.5000 1.1000 0.5000
                 1.1000 1.8700 0.9800 1.8700 0.9800 0.3800 2.0100 0.3800 2.0100 0.3600 2.2500 0.3600
                 2.2500 0.3800 2.4500 0.3800 2.4500 0.8400 2.9300 0.8400 2.9300 0.4400 3.7700 0.4400
                 3.7700 1.2500 4.0700 1.2500 ;
        POLYGON  3.6500 1.7700 3.4100 1.7700 3.4100 1.4400 2.3700 1.4400 2.3700 1.3200 3.1700 1.3200
                 3.1700 0.6800 3.4100 0.6800 3.4100 0.8000 3.2900 0.8000 3.2900 1.3200 3.5300 1.3200
                 3.5300 1.6500 3.6500 1.6500 ;
        POLYGON  3.5300 2.2500 2.9300 2.2500 2.9300 1.9200 2.4500 1.9200 2.4500 2.2500 1.9900 2.2500
                 1.9900 2.1300 2.3300 2.1300 2.3300 1.8000 3.0500 1.8000 3.0500 2.1300 3.5300 2.1300 ;
        POLYGON  3.0300 1.2000 1.9700 1.2000 1.9700 1.7700 1.7300 1.7700 1.7300 1.6500 1.8500 1.6500
                 1.8500 0.6800 2.0900 0.6800 2.0900 0.8000 1.9700 0.8000 1.9700 1.0800 3.0300 1.0800 ;
        POLYGON  0.8400 1.1300 0.7200 1.1300 0.7200 1.0100 0.2400 1.0100 0.2400 1.7200 0.2600 1.7200
                 0.2600 1.9600 0.1400 1.9600 0.1400 1.8400 0.1200 1.8400 0.1200 0.7700 0.1400 0.7700
                 0.1400 0.5300 0.2600 0.5300 0.2600 0.8900 0.8400 0.8900 ;
    END
END EDFFXL

MACRO EDFFX4
    CLASS CORE ;
    FOREIGN EDFFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1600 0.5100 1.6300 ;
        RECT  0.3750 1.1600 0.4950 1.6600 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3650 1.2950 5.6050 1.4900 ;
        RECT  5.2350 1.2300 5.4950 1.4500 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3050 1.2500 6.8950 1.3700 ;
        RECT  6.3950 1.2300 6.6550 1.3800 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.6950 1.3150 8.8150 2.2100 ;
        RECT  7.9000 1.3150 8.8150 1.4350 ;
        RECT  7.4450 0.7200 8.6450 0.8400 ;
        RECT  7.9000 1.1750 8.0500 1.4350 ;
        RECT  7.9000 0.7200 8.0200 1.5550 ;
        RECT  7.8550 1.4350 7.9750 2.2100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3650 0.7200 10.5650 0.8400 ;
        RECT  10.3750 1.3200 10.4950 2.2100 ;
        RECT  9.6400 1.3200 10.4950 1.4400 ;
        RECT  9.6400 1.1750 9.7900 1.4400 ;
        RECT  9.6400 0.7200 9.7600 1.5600 ;
        RECT  9.5350 1.4400 9.6550 2.2100 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  10.9250 -0.1800 11.0450 0.7100 ;
        RECT  9.8450 -0.1800 10.0850 0.3600 ;
        RECT  8.8850 -0.1800 9.1250 0.3600 ;
        RECT  7.9250 -0.1800 8.1650 0.3600 ;
        RECT  6.9650 -0.1800 7.2050 0.3200 ;
        RECT  5.1050 -0.1800 5.2250 0.7900 ;
        RECT  4.2050 0.6100 4.4450 0.7300 ;
        RECT  4.2050 -0.1800 4.3250 0.7300 ;
        RECT  2.5450 0.6100 2.7850 0.7300 ;
        RECT  2.5450 -0.1800 2.6650 0.7300 ;
        RECT  0.5550 -0.1800 0.6750 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  10.7950 1.5800 10.9150 2.7900 ;
        RECT  9.9550 1.5600 10.0750 2.7900 ;
        RECT  9.1150 1.5600 9.2350 2.7900 ;
        RECT  8.2750 1.5600 8.3950 2.7900 ;
        RECT  7.4350 1.7400 7.5550 2.7900 ;
        RECT  5.3250 2.1700 5.5650 2.2900 ;
        RECT  5.3250 2.1700 5.4450 2.7900 ;
        RECT  4.3650 2.1700 4.6050 2.2900 ;
        RECT  4.3650 2.1700 4.4850 2.7900 ;
        RECT  2.5450 1.8100 2.7850 1.9300 ;
        RECT  2.5450 1.8100 2.6650 2.7900 ;
        RECT  0.5550 1.7800 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.4650 0.9000 11.3350 0.9000 11.3350 2.2100 11.2150 2.2100 11.2150 1.4600
                 10.6150 1.4600 10.6150 1.2200 10.7350 1.2200 10.7350 1.3400 11.2150 1.3400
                 11.2150 0.7800 11.3450 0.7800 11.3450 0.6600 11.4650 0.6600 ;
        POLYGON  11.0950 1.2200 10.9750 1.2200 10.9750 0.9500 10.6850 0.9500 10.6850 0.6000
                 8.9250 0.6000 8.9250 1.1600 8.6850 1.1600 8.6850 1.0400 8.8050 1.0400 8.8050 0.6000
                 6.2850 0.6000 6.2850 0.7900 6.1650 0.7900 6.1650 0.4900 5.4900 0.4900 5.4900 1.0300
                 4.9850 1.0300 4.9850 1.6900 5.0850 1.6900 5.0850 1.8100 4.8450 1.8100 4.8450 1.6900
                 4.8650 1.6900 4.8650 1.1700 4.1250 1.1700 4.1250 1.0500 4.6850 1.0500 4.6850 0.6500
                 4.8050 0.6500 4.8050 0.7700 4.9850 0.7700 4.9850 0.9100 5.3700 0.9100 5.3700 0.3700
                 6.2850 0.3700 6.2850 0.4800 10.8050 0.4800 10.8050 0.8300 11.0950 0.8300 ;
        POLYGON  7.6950 1.6200 6.6850 1.6200 6.6850 1.8700 6.5650 1.8700 6.5650 1.5000 7.5750 1.5000
                 7.5750 1.2400 7.6950 1.2400 ;
        POLYGON  7.1350 1.8600 7.0150 1.8600 7.0150 1.9800 6.9250 1.9800 6.9250 2.1100 6.4450 2.1100
                 6.4450 2.2500 5.8850 2.2500 5.8850 2.1300 6.3250 2.1300 6.3250 1.6200 6.0650 1.6200
                 6.0650 1.0500 5.9650 1.0500 5.9650 0.9300 6.4050 0.9300 6.4050 0.7200 6.7350 0.7200
                 6.7350 0.8400 6.5250 0.8400 6.5250 1.0500 6.1850 1.0500 6.1850 1.5000 6.4450 1.5000
                 6.4450 1.9900 6.8050 1.9900 6.8050 1.8600 6.8950 1.8600 6.8950 1.7400 7.1350 1.7400 ;
        POLYGON  6.2050 2.0100 5.4100 2.0100 5.4100 2.0500 4.0850 2.0500 4.0850 2.1100 2.9050 2.1100
                 2.9050 1.6900 2.4250 1.6900 2.4250 2.1100 1.5100 2.1100 1.5100 1.9900 1.4850 1.9900
                 1.4850 1.7500 1.3050 1.7500 1.3050 0.7600 1.3650 0.7600 1.3650 0.6400 1.4850 0.6400
                 1.4850 0.8800 1.4250 0.8800 1.4250 1.6300 1.6050 1.6300 1.6050 1.8700 1.6300 1.8700
                 1.6300 1.9900 2.3050 1.9900 2.3050 1.5700 3.0250 1.5700 3.0250 1.9900 3.9650 1.9900
                 3.9650 1.9300 5.2900 1.9300 5.2900 1.8900 5.7250 1.8900 5.7250 0.7300 5.6850 0.7300
                 5.6850 0.6100 5.9250 0.6100 5.9250 0.7300 5.8450 0.7300 5.8450 1.7400 6.2050 1.7400 ;
        POLYGON  4.7450 1.5500 4.7250 1.5500 4.7250 1.7900 3.7450 1.7900 3.7450 1.8100 3.5050 1.8100
                 3.5050 1.6900 3.5650 1.6900 3.5650 0.6400 3.6850 0.6400 3.6850 1.6700 4.6050 1.6700
                 4.6050 1.4300 4.6250 1.4300 4.6250 1.3100 4.7450 1.3100 ;
        POLYGON  3.9850 1.5500 3.8650 1.5500 3.8650 0.5200 3.0250 0.5200 3.0250 0.9700 2.3050 0.9700
                 2.3050 0.5200 1.7250 0.5200 1.7250 1.3700 1.7850 1.3700 1.7850 1.4900 1.5450 1.4900
                 1.5450 1.3700 1.6050 1.3700 1.6050 0.5200 1.1950 0.5200 1.1950 0.5600 1.0950 0.5600
                 1.0950 1.9000 0.9750 1.9000 0.9750 0.4400 1.0750 0.4400 1.0750 0.4000 2.0050 0.4000
                 2.0050 0.3600 2.2450 0.3600 2.2450 0.4000 2.4250 0.4000 2.4250 0.8500 2.9050 0.8500
                 2.9050 0.4000 3.3450 0.4000 3.3450 0.3600 3.5850 0.3600 3.5850 0.4000 3.9850 0.4000 ;
        POLYGON  3.2650 1.8700 3.1450 1.8700 3.1450 1.2100 2.3250 1.2100 2.3250 1.0900 3.1450 1.0900
                 3.1450 0.6400 3.2650 0.6400 ;
        POLYGON  3.0050 1.4500 2.0850 1.4500 2.0850 1.7500 2.0250 1.7500 2.0250 1.8700 1.9050 1.8700
                 1.9050 1.6300 1.9650 1.6300 1.9650 0.8200 1.8450 0.8200 1.8450 0.7000 2.0850 0.7000
                 2.0850 1.3300 3.0050 1.3300 ;
        POLYGON  0.8350 1.1600 0.7150 1.1600 0.7150 1.0400 0.2400 1.0400 0.2400 1.7500 0.2550 1.7500
                 0.2550 1.9900 0.1350 1.9900 0.1350 1.8700 0.1200 1.8700 0.1200 0.8000 0.1350 0.8000
                 0.1350 0.5600 0.2550 0.5600 0.2550 0.9200 0.8350 0.9200 ;
    END
END EDFFX4

MACRO EDFFX2
    CLASS CORE ;
    FOREIGN EDFFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.1500 0.8550 1.3800 ;
        RECT  0.6050 1.1200 0.7250 1.5300 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3750 1.0750 6.6150 1.2800 ;
        RECT  6.4500 1.0750 6.6000 1.4700 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9750 1.2300 7.2350 1.3800 ;
        RECT  5.8350 1.8300 7.1500 1.9500 ;
        RECT  7.0300 1.1400 7.1500 1.9500 ;
        RECT  6.9900 1.1400 7.1500 1.3800 ;
        RECT  5.5150 1.9900 5.9550 2.1100 ;
        RECT  5.8350 1.3900 5.9550 2.1100 ;
        RECT  5.7750 0.9200 5.8950 1.5100 ;
        RECT  5.6550 0.9200 5.8950 1.0400 ;
        RECT  5.3950 2.1300 5.6350 2.2500 ;
        RECT  5.5150 1.9900 5.6350 2.2500 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7300 0.9400 8.1050 1.0900 ;
        RECT  7.7300 0.7400 7.8650 1.0900 ;
        RECT  7.7300 0.7400 7.8500 1.6500 ;
        RECT  7.6900 1.5300 7.8100 2.1800 ;
        RECT  7.6250 0.7400 7.8650 0.8600 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5100 0.7400 8.8250 0.8600 ;
        RECT  8.5300 1.5300 8.6500 2.1800 ;
        RECT  8.5100 0.7400 8.6300 1.6500 ;
        RECT  8.4800 0.8850 8.6300 1.1450 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.0650 -0.1800 9.3050 0.3800 ;
        RECT  8.1650 -0.1800 8.2850 0.3800 ;
        RECT  7.1450 -0.1800 7.3850 0.3800 ;
        RECT  6.2350 -0.1800 6.4750 0.3800 ;
        RECT  4.6950 -0.1800 4.8150 0.7300 ;
        RECT  2.8150 -0.1800 3.0550 0.3200 ;
        RECT  0.7050 0.5800 0.9450 0.7000 ;
        RECT  0.7050 -0.1800 0.8250 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  8.9500 1.5300 9.0700 2.7900 ;
        RECT  8.1100 1.5700 8.2300 2.7900 ;
        RECT  7.2700 1.5300 7.3900 2.7900 ;
        RECT  6.2350 2.0700 6.4750 2.1900 ;
        RECT  6.2350 2.0700 6.3550 2.7900 ;
        RECT  4.5750 1.9700 4.8150 2.0900 ;
        RECT  4.5750 1.9700 4.6950 2.7900 ;
        RECT  2.8150 2.2600 3.0550 2.7900 ;
        RECT  0.7650 1.6500 0.8850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.7850 0.8600 9.6650 0.8600 9.6650 1.3100 9.5500 1.3100 9.5500 1.7700 9.4300 1.7700
                 9.4300 1.3100 8.7500 1.3100 8.7500 1.1900 9.5450 1.1900 9.5450 0.7400 9.7850 0.7400 ;
        POLYGON  9.6650 0.5400 9.5450 0.5400 9.5450 0.6200 8.3450 0.6200 8.3450 1.4500 7.9700 1.4500
                 7.9700 1.2100 8.2250 1.2100 8.2250 0.6200 7.5050 0.6200 7.5050 1.0000 7.5250 1.0000
                 7.5250 1.2400 7.3850 1.2400 7.3850 0.6200 5.8950 0.6200 5.8950 0.4800 5.2350 0.4800
                 5.2350 0.9700 5.2150 0.9700 5.2150 1.4900 5.2950 1.4900 5.2950 1.6100 5.0550 1.6100
                 5.0550 1.4900 5.0950 1.4900 5.0950 0.9700 4.6950 0.9700 4.6950 1.1200 4.3750 1.1200
                 4.3750 1.0000 4.5750 1.0000 4.5750 0.8500 5.1150 0.8500 5.1150 0.3600 6.0150 0.3600
                 6.0150 0.5000 9.4250 0.5000 9.4250 0.4200 9.6650 0.4200 ;
        POLYGON  6.9100 1.7100 6.6700 1.7100 6.6700 1.5900 6.7350 1.5900 6.7350 0.9550 6.2550 0.9550
                 6.2550 1.2600 6.0150 1.2600 6.0150 0.8350 6.6650 0.8350 6.6650 0.7400 6.9050 0.7400
                 6.9050 0.8600 6.8550 0.8600 6.8550 1.5900 6.9100 1.5900 ;
        POLYGON  5.7750 0.7200 5.5350 0.7200 5.5350 1.6300 5.7150 1.6300 5.7150 1.8700 5.5950 1.8700
                 5.5950 1.8500 4.3900 1.8500 4.3900 1.9000 1.7350 1.9000 1.7350 1.6600 1.5750 1.6600
                 1.5750 0.8000 1.5150 0.8000 1.5150 0.6800 1.7550 0.6800 1.7550 0.8000 1.6950 0.8000
                 1.6950 1.5400 1.8550 1.5400 1.8550 1.7800 4.2700 1.7800 4.2700 1.7300 5.4150 1.7300
                 5.4150 0.6000 5.7750 0.6000 ;
        POLYGON  4.9750 1.3300 4.9350 1.3300 4.9350 1.5800 4.1150 1.5800 4.1150 1.6600 3.7750 1.6600
                 3.7750 0.6200 3.8950 0.6200 3.8950 1.4600 4.8150 1.4600 4.8150 1.2100 4.8550 1.2100
                 4.8550 1.0900 4.9750 1.0900 ;
        POLYGON  4.2550 1.3400 4.0150 1.3400 4.0150 0.5000 3.5500 0.5000 3.5500 0.5600 1.9950 0.5600
                 1.9950 1.2200 2.0550 1.2200 2.0550 1.3400 1.8150 1.3400 1.8150 1.2200 1.8750 1.2200
                 1.8750 0.5600 1.3250 0.5600 1.3250 1.6500 1.3050 1.6500 1.3050 1.7700 1.1850 1.7700
                 1.1850 1.5300 1.2050 1.5300 1.2050 0.7600 1.1850 0.7600 1.1850 0.4400 2.2550 0.4400
                 2.2550 0.3600 2.4950 0.3600 2.4950 0.4400 3.4300 0.4400 3.4300 0.3800 3.5750 0.3800
                 3.5750 0.3600 3.8150 0.3600 3.8150 0.3800 4.1350 0.3800 4.1350 1.2200 4.2550 1.2200 ;
        RECT  2.2750 2.0200 3.8550 2.1400 ;
        POLYGON  3.5750 1.6600 3.3350 1.6600 3.3350 1.0200 2.7750 1.0200 2.7750 1.2000 2.6550 1.2000
                 2.6550 0.9000 3.2950 0.9000 3.2950 0.6800 3.5350 0.6800 3.5350 0.8000 3.4550 0.8000
                 3.4550 1.5400 3.5750 1.5400 ;
        POLYGON  3.2150 1.4400 2.3350 1.4400 2.3350 1.6600 2.0950 1.6600 2.0950 1.5400 2.2150 1.5400
                 2.2150 0.8000 2.1150 0.8000 2.1150 0.6800 2.3550 0.6800 2.3550 0.8000 2.3350 0.8000
                 2.3350 1.3200 3.0950 1.3200 3.0950 1.1400 3.2150 1.1400 ;
        POLYGON  1.0850 1.0200 0.8450 1.0200 0.8450 1.0000 0.4650 1.0000 0.4650 1.7700 0.3450 1.7700
                 0.3450 0.5200 0.4650 0.5200 0.4650 0.8800 1.0850 0.8800 ;
    END
END EDFFX2

MACRO EDFFX1
    CLASS CORE ;
    FOREIGN EDFFX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        RECT  0.4350 1.1750 0.8000 1.3550 ;
        RECT  0.4350 1.1150 0.5550 1.3550 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1050 1.1300 6.3850 1.3700 ;
        RECT  6.1050 1.1300 6.3650 1.3900 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5450 1.1750 6.8900 1.4350 ;
        RECT  5.5650 1.5100 6.6650 1.6300 ;
        RECT  6.5450 1.1750 6.6650 1.6300 ;
        RECT  5.1850 2.1300 5.7450 2.2500 ;
        RECT  5.6250 1.5100 5.7450 2.2500 ;
        RECT  5.5650 0.9200 5.6850 1.6300 ;
        RECT  5.4450 0.9200 5.6850 1.0400 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3500 0.8850 7.4700 1.9900 ;
        RECT  7.3150 0.6800 7.4350 1.0250 ;
        RECT  7.3200 0.8850 7.4700 1.1450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0250 0.5900 9.1450 2.2100 ;
        RECT  8.7700 1.1750 9.1450 1.4350 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        RECT  8.5450 -0.1800 8.6650 0.5300 ;
        RECT  7.8300 -0.1800 7.9500 0.4000 ;
        RECT  6.0250 0.4100 6.2650 0.5300 ;
        RECT  6.0250 -0.1800 6.1450 0.5300 ;
        RECT  4.4850 -0.1800 4.6050 0.7700 ;
        RECT  2.5850 0.3500 2.8250 0.4700 ;
        RECT  2.7050 -0.1800 2.8250 0.4700 ;
        RECT  0.5950 -0.1800 0.7150 0.6950 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        RECT  8.6050 1.7300 8.7250 2.7900 ;
        RECT  7.7700 1.3600 7.8900 2.7900 ;
        RECT  6.3650 1.7500 6.4850 2.7900 ;
        RECT  4.3650 2.1300 4.6050 2.2500 ;
        RECT  4.3650 2.1300 4.4850 2.7900 ;
        RECT  2.5850 1.9100 2.8250 2.0300 ;
        RECT  2.5850 1.9100 2.7050 2.7900 ;
        RECT  0.5950 1.5550 0.7150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.6500 1.1800 8.3950 1.1800 8.3950 1.3000 8.3700 1.3000 8.3700 1.5800 8.2500 1.5800
                 8.2500 1.1800 8.2750 1.1800 8.2750 0.6800 8.3950 0.6800 8.3950 1.0600 8.6500 1.0600 ;
        POLYGON  7.7100 1.2400 7.5900 1.2400 7.5900 0.4800 6.5050 0.4800 6.5050 0.7700 5.7850 0.7700
                 5.7850 0.4800 5.0250 0.4800 5.0250 0.7700 5.0450 0.7700 5.0450 1.5100 4.9650 1.5100
                 4.9650 1.6500 5.0850 1.6500 5.0850 1.7700 4.8450 1.7700 4.8450 1.5100 4.3650 1.5100
                 4.3650 1.2700 4.4850 1.2700 4.4850 1.3900 4.9250 1.3900 4.9250 0.8900 4.9050 0.8900
                 4.9050 0.3600 5.9050 0.3600 5.9050 0.6500 6.3850 0.6500 6.3850 0.3600 7.7100 0.3600 ;
        POLYGON  7.1300 1.6750 6.9050 1.6750 6.9050 1.8700 6.7850 1.8700 6.7850 1.5550 7.0100 1.5550
                 7.0100 1.0100 5.9850 1.0100 5.9850 1.3900 5.8650 1.3900 5.8650 0.8900 7.0100 0.8900
                 7.0100 0.7200 6.6250 0.7200 6.6250 0.6000 7.1300 0.6000 ;
        POLYGON  5.5650 0.7200 5.3250 0.7200 5.3250 1.7500 5.5050 1.7500 5.5050 2.0100 4.1800 2.0100
                 4.1800 2.1100 2.9450 2.1100 2.9450 1.7900 2.4650 1.7900 2.4650 2.1100 1.5250 2.1100
                 1.5250 1.8700 1.3450 1.8700 1.3450 0.7400 1.4050 0.7400 1.4050 0.6200 1.5250 0.6200
                 1.5250 0.8600 1.4650 0.8600 1.4650 1.7500 1.6450 1.7500 1.6450 1.9900 2.3450 1.9900
                 2.3450 1.6700 3.0650 1.6700 3.0650 1.9900 4.0600 1.9900 4.0600 1.8900 5.2050 1.8900
                 5.2050 0.6000 5.5650 0.6000 ;
        POLYGON  4.8050 1.1300 4.2450 1.1300 4.2450 1.7700 3.9050 1.7700 3.9050 1.8100 3.6650 1.8100
                 3.6650 1.6900 3.7850 1.6900 3.7850 1.6500 4.1250 1.6500 4.1250 1.1300 3.6650 1.1300
                 3.6650 0.6200 3.7850 0.6200 3.7850 1.0100 4.8050 1.0100 ;
        POLYGON  4.0050 1.5300 3.8850 1.5300 3.8850 1.4100 3.4250 1.4100 3.4250 1.3100 3.3450 1.3100
                 3.3450 1.0700 3.4250 1.0700 3.4250 0.5000 3.0650 0.5000 3.0650 0.7100 2.3450 0.7100
                 2.3450 0.5000 1.7650 0.5000 1.7650 1.3700 1.8250 1.3700 1.8250 1.4900 1.5850 1.4900
                 1.5850 1.3700 1.6450 1.3700 1.6450 0.5000 1.1350 0.5000 1.1350 1.6750 1.0150 1.6750
                 1.0150 0.3800 2.0250 0.3800 2.0250 0.3600 2.2650 0.3600 2.2650 0.3800 2.4650 0.3800
                 2.4650 0.5900 2.9450 0.5900 2.9450 0.3800 3.5450 0.3800 3.5450 1.2900 4.0050 1.2900 ;
        POLYGON  3.3050 0.9500 3.2250 0.9500 3.2250 1.4300 3.3050 1.4300 3.3050 1.8700 3.1850 1.8700
                 3.1850 1.5500 2.5050 1.5500 2.5050 1.4900 2.3850 1.4900 2.3850 1.3700 2.6250 1.3700
                 2.6250 1.4300 3.1050 1.4300 3.1050 0.8300 3.1850 0.8300 3.1850 0.6200 3.3050 0.6200 ;
        POLYGON  2.9850 1.2200 2.1250 1.2200 2.1250 1.7500 2.0650 1.7500 2.0650 1.8700 1.9450 1.8700
                 1.9450 1.6300 2.0050 1.6300 2.0050 0.8000 1.8850 0.8000 1.8850 0.6800 2.1250 0.6800
                 2.1250 1.1000 2.9850 1.1000 ;
        POLYGON  0.8950 1.0550 0.7750 1.0550 0.7750 0.9950 0.2950 0.9950 0.2950 1.6750 0.1750 1.6750
                 0.1750 0.4550 0.2950 0.4550 0.2950 0.8750 0.7750 0.8750 0.7750 0.8150 0.8950 0.8150 ;
    END
END EDFFX1

MACRO EDFFTRXL
    CLASS CORE ;
    FOREIGN EDFFTRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9350 1.0200 2.0550 1.3050 ;
        RECT  1.8100 0.8850 1.9600 1.1850 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6100 1.4650 7.7600 1.7250 ;
        RECT  7.6100 1.3300 7.7300 1.7250 ;
        RECT  7.3750 1.3300 7.7300 1.4500 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1650 1.5200 10.4250 1.6700 ;
        RECT  10.1650 1.2900 10.3850 1.6700 ;
        RECT  9.5050 1.2900 10.3850 1.4100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0900 1.1750 11.2900 1.4500 ;
        RECT  11.0550 1.0400 11.2250 1.3000 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 1.5800 ;
        RECT  1.2300 1.1750 1.4850 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  10.9650 -0.1800 11.0850 0.9200 ;
        RECT  9.3450 0.5700 9.5850 0.6900 ;
        RECT  9.3450 -0.1800 9.4650 0.6900 ;
        RECT  8.8150 0.5700 9.0550 0.6900 ;
        RECT  8.8150 -0.1800 8.9350 0.6900 ;
        RECT  7.6950 0.6000 7.9350 0.7200 ;
        RECT  7.8150 -0.1800 7.9350 0.7200 ;
        RECT  6.2850 -0.1800 6.5250 0.3200 ;
        RECT  4.6850 0.6500 4.9250 0.7700 ;
        RECT  4.6850 -0.1800 4.8050 0.7700 ;
        RECT  3.0850 -0.1800 3.2050 0.3800 ;
        RECT  1.8450 -0.1800 1.9650 0.4000 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  11.0250 1.9600 11.1450 2.7900 ;
        RECT  7.6150 2.2300 7.7350 2.7900 ;
        RECT  6.2050 2.1700 6.4450 2.2900 ;
        RECT  6.2050 2.1700 6.3250 2.7900 ;
        RECT  4.5650 2.1700 4.8050 2.2900 ;
        RECT  4.5650 2.1700 4.6850 2.7900 ;
        RECT  2.9250 1.8900 3.2050 2.0100 ;
        RECT  3.0850 1.7500 3.2050 2.0100 ;
        RECT  2.9250 1.8900 3.0450 2.7900 ;
        RECT  1.8450 1.9800 1.9650 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6250 1.8400 10.8800 1.8400 10.8800 1.9100 10.6150 1.9100 10.6150 2.2300
                 9.8450 2.2300 9.8450 2.1100 10.4950 2.1100 10.4950 1.7900 10.7600 1.7900
                 10.7600 1.7200 11.5050 1.7200 11.5050 0.9200 11.3850 0.9200 11.3850 0.6800
                 11.5050 0.6800 11.5050 0.8000 11.6250 0.8000 ;
        POLYGON  10.6650 1.6000 10.5450 1.6000 10.5450 1.1700 8.5950 1.1700 8.5950 1.0500
                 10.5450 1.0500 10.5450 0.6800 10.6650 0.6800 ;
        POLYGON  10.2250 1.9100 9.9250 1.9100 9.9250 1.6700 9.3250 1.6700 9.3250 1.8500 9.2050 1.8500
                 9.2050 1.4100 8.3550 1.4100 8.3550 0.9600 7.4550 0.9600 7.4550 0.4800 6.7650 0.4800
                 6.7650 0.5600 6.0450 0.5600 6.0450 0.5200 5.9250 0.5200 5.9250 0.4000 6.1650 0.4000
                 6.1650 0.4400 6.6450 0.4400 6.6450 0.3600 7.5750 0.3600 7.5750 0.8400 8.1750 0.8400
                 8.1750 0.5400 8.2950 0.5400 8.2950 0.6600 8.4750 0.6600 8.4750 0.8100 9.7800 0.8100
                 9.7800 0.6300 10.0450 0.6300 10.0450 0.5100 10.1650 0.5100 10.1650 0.7500
                 9.9000 0.7500 9.9000 0.9300 8.4750 0.9300 8.4750 1.2900 9.3250 1.2900 9.3250 1.5500
                 10.0450 1.5500 10.0450 1.7900 10.2250 1.7900 ;
        POLYGON  9.8050 1.9100 9.6850 1.9100 9.6850 2.0900 8.4550 2.0900 8.4550 1.8900 8.3350 1.8900
                 8.3350 1.7700 8.5750 1.7700 8.5750 1.9700 9.5650 1.9700 9.5650 1.7900 9.8050 1.7900 ;
        POLYGON  8.9350 1.8300 8.8150 1.8300 8.8150 1.6500 8.0950 1.6500 8.0950 1.8300 7.9750 1.8300
                 7.9750 1.5300 8.9350 1.5300 ;
        POLYGON  8.2950 2.2100 8.0550 2.2100 8.0550 2.0700 6.7300 2.0700 6.7300 2.0500 6.0550 2.0500
                 6.0550 2.1100 4.9250 2.1100 4.9250 2.0500 4.2500 2.0500 4.2500 2.1100 3.4450 2.1100
                 3.4450 2.2500 3.1650 2.2500 3.1650 2.1300 3.3250 2.1300 3.3250 1.6300 2.9150 1.6300
                 2.9150 1.7700 2.7850 1.7700 2.7850 1.8700 2.6650 1.8700 2.6650 1.8600 1.6850 1.8600
                 1.6850 1.9600 1.4450 1.9600 1.4450 1.8400 1.5650 1.8400 1.5650 1.7400 2.6250 1.7400
                 2.6250 0.9000 2.6050 0.9000 2.6050 0.6600 2.7250 0.6600 2.7250 0.7800 2.7450 0.7800
                 2.7450 1.5100 3.4450 1.5100 3.4450 1.9900 4.1300 1.9900 4.1300 1.9300 5.0450 1.9300
                 5.0450 1.9900 5.9350 1.9900 5.9350 1.9300 6.8500 1.9300 6.8500 1.9500 8.1750 1.9500
                 8.1750 2.0900 8.2950 2.0900 ;
        POLYGON  7.9750 1.2000 7.2550 1.2000 7.2550 1.8300 7.1350 1.8300 7.1350 0.7200 7.0950 0.7200
                 7.0950 0.6000 7.3350 0.6000 7.3350 0.7200 7.2550 0.7200 7.2550 1.0800 7.9750 1.0800 ;
        POLYGON  6.9450 0.8400 6.8850 0.8400 6.8850 1.6900 6.9250 1.6900 6.9250 1.8100 6.6850 1.8100
                 6.6850 1.6900 6.7650 1.6900 6.7650 1.4800 5.6450 1.4800 5.6450 1.3600 6.7650 1.3600
                 6.7650 0.8400 6.7050 0.8400 6.7050 0.7200 6.9450 0.7200 ;
        POLYGON  6.6450 1.1600 5.6850 1.1600 5.6850 0.5400 5.2850 0.5400 5.2850 1.5300 5.1650 1.5300
                 5.1650 1.0100 4.4450 1.0100 4.4450 0.5400 4.0850 0.5400 4.0850 1.5500 3.9650 1.5500
                 3.9650 0.5400 3.4450 0.5400 3.4450 0.6200 2.8450 0.6200 2.8450 0.5400 2.4350 0.5400
                 2.4350 0.6800 2.3350 0.6800 2.3350 0.8000 2.3950 0.8000 2.3950 1.5800 2.2750 1.5800
                 2.2750 0.9200 2.2150 0.9200 2.2150 0.5600 2.3150 0.5600 2.3150 0.4200 2.9650 0.4200
                 2.9650 0.5000 3.3250 0.5000 3.3250 0.4200 3.4450 0.4200 3.4450 0.3800 3.6850 0.3800
                 3.6850 0.4200 4.5650 0.4200 4.5650 0.8900 5.1650 0.8900 5.1650 0.4200 5.8050 0.4200
                 5.8050 1.0400 6.6450 1.0400 ;
        POLYGON  5.5650 1.2400 5.5250 1.2400 5.5250 1.8700 5.4050 1.8700 5.4050 1.7700 4.9250 1.7700
                 4.9250 1.4900 4.4450 1.4900 4.4450 1.3700 5.0450 1.3700 5.0450 1.6500 5.4050 1.6500
                 5.4050 1.1200 5.4450 1.1200 5.4450 0.6600 5.5650 0.6600 ;
        POLYGON  5.0250 1.2500 4.3250 1.2500 4.3250 1.8100 4.0850 1.8100 4.0850 1.6900 4.2050 1.6900
                 4.2050 0.6600 4.3250 0.6600 4.3250 1.1300 5.0250 1.1300 ;
        POLYGON  3.8450 1.8700 3.7250 1.8700 3.7250 1.3900 2.8650 1.3900 2.8650 1.2700 3.7250 1.2700
                 3.7250 0.8400 3.6050 0.8400 3.6050 0.7200 3.8450 0.7200 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END EDFFTRXL

MACRO EDFFTRX4
    CLASS CORE ;
    FOREIGN EDFFTRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 15.0800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1750 0.6450 1.4100 ;
        RECT  0.5250 1.1700 0.6450 1.4100 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0150 1.2500 2.3950 1.3700 ;
        RECT  1.0250 1.8100 2.1350 1.9300 ;
        RECT  2.0150 1.2500 2.1350 1.9300 ;
        RECT  1.0250 1.1700 1.1450 1.9300 ;
        RECT  0.8850 1.5200 1.1450 1.6700 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6550 1.2300 5.0350 1.4200 ;
        RECT  4.6550 1.2300 4.9150 1.4450 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 1.2200 9.5550 1.4500 ;
        RECT  9.3050 1.0400 9.4250 1.4500 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.8850 1.4900 12.1250 1.6100 ;
        RECT  11.3250 0.8500 12.1050 0.9700 ;
        RECT  11.9850 0.6800 12.1050 0.9700 ;
        RECT  11.3250 1.3700 12.0050 1.4900 ;
        RECT  11.3250 1.1750 11.5300 1.4900 ;
        RECT  10.9250 1.4900 11.4450 1.6100 ;
        RECT  11.3250 0.8000 11.4450 1.6100 ;
        RECT  11.1450 0.8000 11.4450 0.9200 ;
        RECT  11.1450 0.6800 11.2650 0.9200 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.8050 1.4900 14.0450 1.6100 ;
        RECT  12.8450 1.3800 13.9250 1.5000 ;
        RECT  12.8600 0.8500 13.7850 0.9700 ;
        RECT  13.6650 0.6800 13.7850 0.9700 ;
        RECT  12.8450 1.3800 13.0850 1.6100 ;
        RECT  12.8300 1.1750 12.9800 1.4350 ;
        RECT  12.8600 0.8000 12.9800 1.6100 ;
        RECT  12.8250 0.6800 12.9450 0.9200 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 15.0800 0.1800 ;
        RECT  14.0850 -0.1800 14.2050 0.7300 ;
        RECT  13.2450 -0.1800 13.3650 0.7300 ;
        RECT  12.4050 -0.1800 12.5250 0.7300 ;
        RECT  11.5650 -0.1800 11.6850 0.7300 ;
        RECT  10.7250 -0.1800 10.8450 0.7300 ;
        RECT  9.8250 -0.1800 9.9450 0.8200 ;
        RECT  8.1750 0.7000 8.4150 0.8200 ;
        RECT  8.1750 -0.1800 8.2950 0.8200 ;
        RECT  6.4550 0.5300 6.6950 0.6500 ;
        RECT  6.4550 -0.1800 6.5750 0.6500 ;
        RECT  4.7350 -0.1800 4.9750 0.3400 ;
        RECT  3.7750 -0.1800 3.8950 0.3800 ;
        RECT  2.6450 0.5300 2.8850 0.6500 ;
        RECT  2.6450 -0.1800 2.7650 0.6500 ;
        RECT  2.2550 0.5300 2.4950 0.6500 ;
        RECT  2.3750 -0.1800 2.4950 0.6500 ;
        RECT  0.8050 -0.1800 0.9250 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 15.0800 2.7900 ;
        RECT  14.2850 1.9700 14.5250 2.0900 ;
        RECT  14.2850 1.9700 14.4050 2.7900 ;
        RECT  13.3250 1.9700 13.5650 2.0900 ;
        RECT  13.3250 1.9700 13.4450 2.7900 ;
        RECT  12.3650 1.9700 12.6050 2.0900 ;
        RECT  12.3650 1.9700 12.4850 2.7900 ;
        RECT  11.4050 1.9700 11.6450 2.0900 ;
        RECT  11.4050 1.9700 11.5250 2.7900 ;
        RECT  10.4450 1.9700 10.6850 2.0900 ;
        RECT  10.4450 1.9700 10.5650 2.7900 ;
        RECT  9.5650 2.2900 9.8050 2.7900 ;
        RECT  8.3350 2.2900 8.5750 2.7900 ;
        RECT  6.5550 2.1100 6.6750 2.7900 ;
        RECT  5.2550 2.1500 5.3750 2.7900 ;
        RECT  4.4450 2.1700 4.5650 2.7900 ;
        RECT  0.7850 2.2900 1.0250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  14.9450 2.0800 14.8250 2.0800 14.8250 1.5500 14.5850 1.5500 14.5850 0.9700
                 14.0450 0.9700 14.0450 1.2600 13.9250 1.2600 13.9250 0.8500 14.5050 0.8500
                 14.5050 0.6800 14.6250 0.6800 14.6250 0.8000 14.7050 0.8000 14.7050 1.4300
                 14.9450 1.4300 ;
        POLYGON  14.4650 1.8500 10.1450 1.8500 10.1450 1.9500 10.0400 1.9500 10.0400 2.1700
                 8.0650 2.1700 8.0650 2.1500 7.0050 2.1500 7.0050 1.9900 6.3300 1.9900 6.3300 2.0300
                 5.0050 2.0300 5.0050 2.0500 3.9450 2.0500 3.9450 2.2500 3.8250 2.2500 3.8250 1.9300
                 4.8850 1.9300 4.8850 1.9100 6.2100 1.9100 6.2100 1.8700 7.1250 1.8700 7.1250 2.0300
                 8.2550 2.0300 8.2550 2.0500 9.9200 2.0500 9.9200 1.8300 10.0250 1.8300 10.0250 1.4300
                 10.2450 1.4300 10.2450 0.6800 10.3650 0.6800 10.3650 1.1700 11.0450 1.1700
                 11.0450 1.2900 10.3650 1.2900 10.3650 1.5500 10.1450 1.5500 10.1450 1.7300
                 14.3450 1.7300 14.3450 1.0900 14.4650 1.0900 ;
        POLYGON  10.1050 1.3100 9.9050 1.3100 9.9050 1.7100 9.6400 1.7100 9.6400 1.9300 8.3750 1.9300
                 8.3750 1.9100 7.4550 1.9100 7.4550 1.5500 7.5350 1.5500 7.5350 0.6400 7.6550 0.6400
                 7.6550 1.6700 7.5750 1.6700 7.5750 1.7900 8.4950 1.7900 8.4950 1.8100 9.5200 1.8100
                 9.5200 1.5900 9.7850 1.5900 9.7850 1.1900 9.9850 1.1900 9.9850 1.0700 10.1050 1.0700 ;
        POLYGON  9.4650 0.9200 9.1750 0.9200 9.1750 1.5700 9.3250 1.5700 9.3250 1.6900 9.0550 1.6900
                 9.0550 0.8000 9.3450 0.8000 9.3450 0.6800 9.0800 0.6800 9.0800 0.5200 8.6550 0.5200
                 8.6550 1.0600 7.9350 1.0600 7.9350 0.5200 7.4150 0.5200 7.4150 1.4300 7.2950 1.4300
                 7.2950 0.5200 6.9350 0.5200 6.9350 0.8900 6.0550 0.8900 6.0550 1.4300 5.9350 1.4300
                 5.9350 0.4800 5.4550 0.4800 5.4550 0.3600 6.0550 0.3600 6.0550 0.7700 6.8150 0.7700
                 6.8150 0.4000 7.6950 0.4000 7.6950 0.3600 7.9350 0.3600 7.9350 0.4000 8.0550 0.4000
                 8.0550 0.9400 8.5350 0.9400 8.5350 0.4800 8.4350 0.4800 8.4350 0.3600 8.6750 0.3600
                 8.6750 0.4000 9.2000 0.4000 9.2000 0.5600 9.4650 0.5600 ;
        POLYGON  8.9350 1.6900 8.6950 1.6900 8.6950 1.5700 8.7750 1.5700 8.7750 1.3700 7.7750 1.3700
                 7.7750 1.2500 8.7750 1.2500 8.7750 0.6400 8.8950 0.6400 8.8950 1.5700 8.9350 1.5700 ;
        POLYGON  7.1750 1.4900 7.1550 1.4900 7.1550 1.7500 7.0350 1.7500 7.0350 1.4900 6.5750 1.4900
                 6.5750 1.3700 6.4150 1.3700 6.4150 1.2500 6.6950 1.2500 6.6950 1.3700 7.0550 1.3700
                 7.0550 0.6400 7.1750 0.6400 ;
        POLYGON  6.9350 1.2500 6.8150 1.2500 6.8150 1.1300 6.2950 1.1300 6.2950 1.6700 6.0350 1.6700
                 6.0350 1.6900 5.6950 1.6900 5.6950 0.8200 5.5750 0.8200 5.5750 0.7000 5.8150 0.7000
                 5.8150 1.5500 6.1750 1.5500 6.1750 1.0100 6.9350 1.0100 ;
        POLYGON  5.3350 0.4800 5.2150 0.4800 5.2150 0.5800 4.1350 0.5800 4.1350 0.6600 3.6850 0.6600
                 3.6850 1.1300 2.8550 1.1300 2.8550 1.7500 2.7350 1.7500 2.7350 1.1300 1.8250 1.1300
                 1.8250 1.5700 1.8950 1.5700 1.8950 1.6900 1.6550 1.6900 1.6550 1.5700 1.7050 1.5700
                 1.7050 0.7200 1.5550 0.7200 1.5550 0.6000 1.8250 0.6000 1.8250 1.0100 3.5650 1.0100
                 3.5650 0.5400 4.0150 0.5400 4.0150 0.4600 5.0950 0.4600 5.0950 0.3600 5.3350 0.3600 ;
        POLYGON  4.9550 1.6900 4.3750 1.6900 4.3750 1.2300 4.1750 1.2300 4.1750 1.1100 4.3750 1.1100
                 4.3750 0.8200 4.2550 0.8200 4.2550 0.7000 4.4950 0.7000 4.4950 1.5700 4.9550 1.5700 ;
        POLYGON  4.0850 1.8100 3.9650 1.8100 3.9650 1.5700 3.2450 1.5700 3.2450 1.8100 3.1250 1.8100
                 3.1250 1.4500 4.0850 1.4500 ;
        POLYGON  3.6650 2.0500 2.3750 2.0500 2.3750 1.8100 2.2550 1.8100 2.2550 1.6900 2.4950 1.6900
                 2.4950 1.9300 3.5450 1.9300 3.5450 1.6900 3.6650 1.6900 ;
        POLYGON  3.2450 0.5200 3.1250 0.5200 3.1250 0.8900 1.9450 0.8900 1.9450 0.4800 1.3450 0.4800
                 1.3450 0.8000 1.3850 0.8000 1.3850 1.5700 1.5050 1.5700 1.5050 1.6900 1.2650 1.6900
                 1.2650 0.9200 1.2250 0.9200 1.2250 0.3600 2.0650 0.3600 2.0650 0.7700 3.0050 0.7700
                 3.0050 0.4000 3.2450 0.4000 ;
        POLYGON  2.0550 2.1700 0.3650 2.1700 0.3650 1.6750 0.1200 1.6750 0.1200 0.9300 0.3850 0.9300
                 0.3850 0.6800 0.5050 0.6800 0.5050 1.0500 0.2400 1.0500 0.2400 1.5550 0.4850 1.5550
                 0.4850 2.0500 2.0550 2.0500 ;
    END
END EDFFTRX4

MACRO EDFFTRX2
    CLASS CORE ;
    FOREIGN EDFFTRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.3400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1750 0.6450 1.4100 ;
        RECT  0.5250 1.1700 0.6450 1.4100 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0150 1.2500 2.4050 1.3700 ;
        RECT  1.0250 1.8100 2.1350 1.9300 ;
        RECT  2.0150 1.2500 2.1350 1.9300 ;
        RECT  1.0250 1.1700 1.1450 1.9300 ;
        RECT  0.8850 1.5200 1.1450 1.6700 ;
        END
    END E
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4650 1.2500 4.5850 1.5600 ;
        RECT  4.4200 1.4400 4.5700 1.7550 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.2300 10.7150 1.4450 ;
        RECT  10.5650 0.9700 10.6850 1.4450 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.2550 1.1750 11.5300 1.4350 ;
        RECT  11.1150 1.5500 11.3750 1.6700 ;
        RECT  11.2550 0.5900 11.3750 1.6700 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  12.0750 1.5500 12.3150 1.6700 ;
        RECT  12.0750 1.1750 12.2150 1.6700 ;
        RECT  12.0950 0.5900 12.2150 1.6700 ;
        RECT  11.9600 1.1750 12.2150 1.4350 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.3400 0.1800 ;
        RECT  12.5150 -0.1800 12.6350 0.6400 ;
        RECT  11.6750 -0.1800 11.7950 0.6400 ;
        RECT  10.8350 -0.1800 10.9550 0.7900 ;
        RECT  9.4850 -0.1800 9.7250 0.3800 ;
        RECT  7.5850 0.5300 7.8250 0.6500 ;
        RECT  7.5850 -0.1800 7.7050 0.6500 ;
        RECT  5.5650 0.5300 5.8050 0.6500 ;
        RECT  5.6850 -0.1800 5.8050 0.6500 ;
        RECT  4.1550 -0.1800 4.2750 0.6500 ;
        RECT  2.7550 0.5300 2.9950 0.6500 ;
        RECT  2.7550 -0.1800 2.8750 0.6500 ;
        RECT  2.4250 -0.1800 2.5450 0.6500 ;
        RECT  0.8450 -0.1800 0.9650 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.3400 2.7900 ;
        RECT  12.6150 2.1500 12.7350 2.7900 ;
        RECT  11.5950 2.0300 11.8350 2.1500 ;
        RECT  11.5950 2.0300 11.7150 2.7900 ;
        RECT  10.6950 2.0900 10.8150 2.7900 ;
        RECT  9.4250 1.6800 9.6650 1.8100 ;
        RECT  9.4250 1.6800 9.5450 2.7900 ;
        RECT  7.5850 2.2900 7.8250 2.7900 ;
        RECT  5.6250 2.1500 5.7450 2.7900 ;
        RECT  4.4450 2.2100 4.5650 2.7900 ;
        RECT  0.7850 2.2900 1.0250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.2050 1.7300 13.0850 1.7300 13.0850 1.3500 12.3350 1.3500 12.3350 1.2300
                 12.9950 1.2300 12.9950 0.5900 13.1150 0.5900 13.1150 1.2300 13.2050 1.2300 ;
        POLYGON  13.0550 2.1900 12.9350 2.1900 12.9350 2.0300 12.7300 2.0300 12.7300 1.9100
                 10.8200 1.9100 10.8200 1.9700 10.0250 1.9700 10.0250 2.1600 9.9050 2.1600
                 9.9050 1.5600 9.3050 1.5600 9.3050 2.2100 9.1850 2.2100 9.1850 2.1700 6.2100 2.1700
                 6.2100 2.0300 5.2700 2.0300 5.2700 2.0500 5.0050 2.0500 5.0050 2.0900 3.9450 2.0900
                 3.9450 2.2500 3.8250 2.2500 3.8250 1.9700 4.8850 1.9700 4.8850 1.9300 5.1500 1.9300
                 5.1500 1.9100 6.3300 1.9100 6.3300 2.0500 9.1650 2.0500 9.1650 1.4400 9.9050 1.4400
                 9.9050 0.7400 10.2050 0.7400 10.2050 0.8600 10.0250 0.8600 10.0250 1.8500
                 10.7000 1.8500 10.7000 1.7900 10.8750 1.7900 10.8750 1.2900 10.9750 1.2900
                 10.9750 0.9100 11.0950 0.9100 11.0950 1.4100 10.9950 1.4100 10.9950 1.7900
                 12.8500 1.7900 12.8500 1.9100 13.0550 1.9100 ;
        POLYGON  10.5350 0.7900 10.4450 0.7900 10.4450 1.1100 10.3350 1.1100 10.3350 1.7300
                 10.2150 1.7300 10.2150 0.9900 10.3250 0.9900 10.3250 0.6200 9.1900 0.6200
                 9.1900 0.5000 8.5450 0.5000 8.5450 1.2500 8.5650 1.2500 8.5650 1.3700 8.3250 1.3700
                 8.3250 1.2500 8.4250 1.2500 8.4250 0.5000 8.0650 0.5000 8.0650 0.8900 7.2050 0.8900
                 7.2050 1.4300 7.0850 1.4300 7.0850 0.5600 6.4050 0.5600 6.4050 1.1300 5.4150 1.1300
                 5.4150 1.0100 6.2850 1.0100 6.2850 0.4400 7.2050 0.4400 7.2050 0.7700 7.9450 0.7700
                 7.9450 0.3800 8.9250 0.3800 8.9250 0.3600 9.1650 0.3600 9.1650 0.3800 9.3100 0.3800
                 9.3100 0.5000 10.5350 0.5000 ;
        POLYGON  9.7450 1.2400 9.6250 1.2400 9.6250 1.0800 8.8050 1.0800 8.8050 1.6900 8.5650 1.6900
                 8.5650 1.5700 8.6850 1.5700 8.6850 0.8400 8.8450 0.8400 8.8450 0.6200 8.9650 0.6200
                 8.9650 0.9600 9.7450 0.9600 ;
        POLYGON  9.1650 1.3200 9.0450 1.3200 9.0450 1.9300 6.5400 1.9300 6.5400 1.4900 6.4850 1.4900
                 6.4850 1.3700 5.3150 1.3700 5.3150 1.7500 5.1950 1.7500 5.1950 1.4900 5.1750 1.4900
                 5.1750 1.1300 4.9650 1.1300 4.9650 0.6800 5.2050 0.6800 5.2050 1.0100 5.2950 1.0100
                 5.2950 1.2500 6.7250 1.2500 6.7250 1.3700 6.6600 1.3700 6.6600 1.8100 8.9250 1.8100
                 8.9250 1.2000 9.1650 1.2000 ;
        POLYGON  8.3050 1.1300 8.2050 1.1300 8.2050 1.5700 8.3050 1.5700 8.3050 1.6900 8.0650 1.6900
                 8.0650 1.5700 8.0850 1.5700 8.0850 1.1300 7.6050 1.1300 7.6050 1.1400 7.3650 1.1400
                 7.3650 1.0200 7.4850 1.0200 7.4850 1.0100 8.1850 1.0100 8.1850 0.6200 8.3050 0.6200 ;
        POLYGON  7.9650 1.3700 7.8450 1.3700 7.8450 1.6700 7.0200 1.6700 7.0200 1.6900 6.7800 1.6900
                 6.7800 1.5700 6.8450 1.5700 6.8450 0.8000 6.5250 0.8000 6.5250 0.6800 6.9650 0.6800
                 6.9650 1.5500 7.7250 1.5500 7.7250 1.2500 7.9650 1.2500 ;
        POLYGON  6.1650 0.4800 6.0450 0.4800 6.0450 0.8900 5.3250 0.8900 5.3250 0.5600 5.1900 0.5600
                 5.1900 0.5000 4.5150 0.5000 4.5150 0.8900 3.7950 0.8900 3.7950 1.1300 2.8550 1.1300
                 2.8550 1.7500 2.7350 1.7500 2.7350 1.1300 1.8950 1.1300 1.8950 1.6900 1.6550 1.6900
                 1.6550 1.5700 1.7750 1.5700 1.7750 1.0100 1.7250 1.0100 1.7250 0.6000 1.8450 0.6000
                 1.8450 0.8900 1.8950 0.8900 1.8950 1.0100 3.6750 1.0100 3.6750 0.6200 3.7950 0.6200
                 3.7950 0.7400 3.9850 0.7400 3.9850 0.7700 4.3950 0.7700 4.3950 0.3800 5.3100 0.3800
                 5.3100 0.4400 5.4450 0.4400 5.4450 0.7700 5.9250 0.7700 5.9250 0.3600 6.1650 0.3600 ;
        POLYGON  4.9250 1.8100 4.8050 1.8100 4.8050 1.6900 4.7050 1.6900 4.7050 1.1300 4.2450 1.1300
                 4.2450 1.2500 4.1250 1.2500 4.1250 1.0100 4.6350 1.0100 4.6350 0.6200 4.7550 0.6200
                 4.7550 0.8900 4.8250 0.8900 4.8250 1.5700 4.9250 1.5700 ;
        POLYGON  4.0850 1.8100 3.9650 1.8100 3.9650 1.5700 3.2450 1.5700 3.2450 1.8100 3.1250 1.8100
                 3.1250 1.4500 4.0850 1.4500 ;
        POLYGON  3.6650 2.0500 2.3750 2.0500 2.3750 1.8100 2.2550 1.8100 2.2550 1.6900 2.4950 1.6900
                 2.4950 1.9300 3.5450 1.9300 3.5450 1.6900 3.6650 1.6900 ;
        POLYGON  3.3550 0.4800 3.2350 0.4800 3.2350 0.8900 2.0550 0.8900 2.0550 0.4800 1.3850 0.4800
                 1.3850 1.5700 1.5050 1.5700 1.5050 1.6900 1.2650 1.6900 1.2650 0.3600 2.1750 0.3600
                 2.1750 0.7700 3.1150 0.7700 3.1150 0.3600 3.3550 0.3600 ;
        POLYGON  2.0650 2.1700 0.3650 2.1700 0.3650 1.6750 0.1200 1.6750 0.1200 0.9300 0.4250 0.9300
                 0.4250 0.6800 0.5450 0.6800 0.5450 1.0500 0.2400 1.0500 0.2400 1.5550 0.4850 1.5550
                 0.4850 2.0500 2.0650 2.0500 ;
    END
END EDFFTRX2

MACRO EDFFTRX1
    CLASS CORE ;
    FOREIGN EDFFTRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9450 1.1000 2.0800 1.3400 ;
        RECT  1.8100 1.1750 1.9750 1.4350 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5600 1.3500 7.8000 1.5200 ;
        RECT  7.6100 1.3500 7.7600 1.7250 ;
        END
    END RN
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.5200 10.7150 1.6700 ;
        RECT  10.4550 1.3200 10.6750 1.6700 ;
        RECT  9.7950 1.3200 10.6750 1.4400 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.3300 1.1750 11.5300 1.4500 ;
        RECT  11.3450 1.0400 11.5150 1.4500 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2888  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3800 0.6800 1.5000 1.0250 ;
        RECT  1.3300 0.8850 1.4500 2.2100 ;
        RECT  1.2300 0.8850 1.4500 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.2550 -0.1800 11.3750 0.9200 ;
        RECT  9.5350 0.6000 9.7750 0.7200 ;
        RECT  9.5350 -0.1800 9.6550 0.7200 ;
        RECT  8.9400 0.6000 9.1800 0.7200 ;
        RECT  8.9400 -0.1800 9.0600 0.7200 ;
        RECT  7.8800 0.6000 8.1200 0.7200 ;
        RECT  8.0000 -0.1800 8.1200 0.7200 ;
        RECT  6.4100 -0.1800 6.6500 0.3200 ;
        RECT  4.8100 0.5700 5.0500 0.6900 ;
        RECT  4.8100 -0.1800 4.9300 0.6900 ;
        RECT  3.0900 0.6800 3.3300 0.8000 ;
        RECT  3.2100 -0.1800 3.3300 0.8000 ;
        RECT  1.8000 -0.1800 1.9200 0.9200 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.3150 1.9600 11.4350 2.7900 ;
        RECT  7.7850 2.2200 7.9050 2.7900 ;
        RECT  6.3100 2.1700 6.5500 2.2900 ;
        RECT  6.3100 2.1700 6.4300 2.7900 ;
        RECT  4.7100 2.2300 4.8300 2.7900 ;
        RECT  3.0100 1.8700 3.2700 1.9900 ;
        RECT  3.1500 1.6400 3.2700 1.9900 ;
        RECT  3.0100 1.8700 3.1300 2.7900 ;
        RECT  1.7500 2.1000 1.9900 2.2200 ;
        RECT  1.7500 2.1000 1.8700 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.9150 1.8400 11.1200 1.8400 11.1200 2.1500 10.3750 2.1500 10.3750 2.2400
                 10.1350 2.2400 10.1350 2.1200 10.2550 2.1200 10.2550 2.0300 11.0000 2.0300
                 11.0000 1.7200 11.7950 1.7200 11.7950 0.9200 11.6750 0.9200 11.6750 0.6800
                 11.7950 0.6800 11.7950 0.8000 11.9150 0.8000 ;
        POLYGON  10.9550 1.6000 10.8350 1.6000 10.8350 1.2000 8.8850 1.2000 8.8850 1.0800
                 10.8350 1.0800 10.8350 0.6800 10.9550 0.6800 ;
        POLYGON  10.5150 1.9100 10.2150 1.9100 10.2150 1.6800 9.6150 1.6800 9.6150 1.8600 9.4950 1.8600
                 9.4950 1.4400 8.6450 1.4400 8.6450 0.9600 7.6400 0.9600 7.6400 0.4800 6.8900 0.4800
                 6.8900 0.5600 6.1700 0.5600 6.1700 0.4800 6.0500 0.4800 6.0500 0.3600 6.2900 0.3600
                 6.2900 0.4400 6.7700 0.4400 6.7700 0.3600 7.7600 0.3600 7.7600 0.8400 8.3600 0.8400
                 8.3600 0.5400 8.4800 0.5400 8.4800 0.6600 8.7650 0.6600 8.7650 0.8400 9.9100 0.8400
                 9.9100 0.6000 10.4150 0.6000 10.4150 0.7200 10.0300 0.7200 10.0300 0.9600
                 8.7650 0.9600 8.7650 1.3200 9.6150 1.3200 9.6150 1.5600 10.3350 1.5600 10.3350 1.7900
                 10.5150 1.7900 ;
        POLYGON  10.0950 1.9200 9.9750 1.9200 9.9750 2.1000 8.7450 2.1000 8.7450 1.9200 8.6250 1.9200
                 8.6250 1.8000 8.8650 1.8000 8.8650 1.9800 9.8550 1.9800 9.8550 1.8000 10.0950 1.8000 ;
        POLYGON  9.2250 1.8600 9.1050 1.8600 9.1050 1.6800 8.3850 1.6800 8.3850 1.8600 8.2650 1.8600
                 8.2650 1.5600 9.2250 1.5600 ;
        POLYGON  8.5850 2.2400 8.3450 2.2400 8.3450 2.1000 7.0200 2.1000 7.0200 2.0500 6.1900 2.0500
                 6.1900 2.1100 3.5100 2.1100 3.5100 2.2500 3.2500 2.2500 3.2500 2.1300 3.3900 2.1300
                 3.3900 1.5200 2.8500 1.5200 2.8500 1.9900 2.7300 1.9900 2.7300 1.9800 1.5700 1.9800
                 1.5700 1.2400 1.6900 1.2400 1.6900 1.8600 2.6300 1.8600 2.6300 1.5900 2.6100 1.5900
                 2.6100 0.6800 2.7300 0.6800 2.7300 1.4000 3.5100 1.4000 3.5100 1.9900 6.0700 1.9900
                 6.0700 1.9300 7.1400 1.9300 7.1400 1.9800 8.4650 1.9800 8.4650 2.1200 8.5850 2.1200 ;
        POLYGON  8.1650 1.2300 7.4400 1.2300 7.4400 1.7400 7.4250 1.7400 7.4250 1.8600 7.3050 1.8600
                 7.3050 1.6200 7.3200 1.6200 7.3200 0.7200 7.2800 0.7200 7.2800 0.6000 7.5200 0.6000
                 7.5200 0.7200 7.4400 0.7200 7.4400 1.1100 8.1650 1.1100 ;
        POLYGON  7.1300 0.8000 7.0100 0.8000 7.0100 1.6900 7.0300 1.6900 7.0300 1.8100 6.7900 1.8100
                 6.7900 1.6900 6.8900 1.6900 6.8900 1.4400 5.7500 1.4400 5.7500 1.3200 6.8900 1.3200
                 6.8900 0.6800 7.1300 0.6800 ;
        POLYGON  6.7500 1.1200 5.7900 1.1200 5.7900 1.0000 5.8100 1.0000 5.8100 0.5000 5.3900 0.5000
                 5.3900 1.5500 5.2700 1.5500 5.2700 0.9300 4.5700 0.9300 4.5700 0.5000 4.2100 0.5000
                 4.2100 1.3700 4.2700 1.3700 4.2700 1.4900 4.0300 1.4900 4.0300 1.3700 4.0900 1.3700
                 4.0900 0.5000 3.5700 0.5000 3.5700 1.0400 2.8500 1.0400 2.8500 0.5600 2.3400 0.5600
                 2.3400 0.8000 2.3500 0.8000 2.3500 1.6200 2.4700 1.6200 2.4700 1.7400 2.2300 1.7400
                 2.2300 0.9200 2.2200 0.9200 2.2200 0.4400 2.9700 0.4400 2.9700 0.9200 3.4500 0.9200
                 3.4500 0.3800 3.5900 0.3800 3.5900 0.3600 3.8300 0.3600 3.8300 0.3800 4.6900 0.3800
                 4.6900 0.8100 5.2700 0.8100 5.2700 0.3800 5.9300 0.3800 5.9300 1.0000 6.7500 1.0000 ;
        POLYGON  5.6900 0.8600 5.6300 0.8600 5.6300 1.8700 5.5100 1.8700 5.5100 1.7900 5.0300 1.7900
                 5.0300 1.4900 4.6300 1.4900 4.6300 1.3700 5.1500 1.3700 5.1500 1.6700 5.5100 1.6700
                 5.5100 0.7400 5.5700 0.7400 5.5700 0.6200 5.6900 0.6200 ;
        POLYGON  5.0900 1.1700 4.5100 1.1700 4.5100 1.7300 4.3500 1.7300 4.3500 1.8700 4.2300 1.8700
                 4.2300 1.6100 4.3900 1.6100 4.3900 1.1700 4.3300 1.1700 4.3300 0.6200 4.4500 0.6200
                 4.4500 1.0500 5.0900 1.0500 ;
        POLYGON  3.9700 0.8000 3.9100 0.8000 3.9100 1.6300 3.9300 1.6300 3.9300 1.8700 3.8100 1.8700
                 3.8100 1.7500 3.7900 1.7500 3.7900 1.2800 2.9500 1.2800 2.9500 1.1600 3.7900 1.1600
                 3.7900 0.8000 3.7300 0.8000 3.7300 0.6800 3.9700 0.6800 ;
        POLYGON  1.1400 1.5800 1.0200 1.5800 1.0200 1.3850 0.9900 1.3850 0.9900 1.2000 0.3750 1.2000
                 0.3750 1.0800 0.9900 1.0800 0.9900 0.6800 1.1100 0.6800 1.1100 1.2650 1.1400 1.2650 ;
    END
END EDFFTRX1

MACRO EDFFHQX8
    CLASS CORE ;
    FOREIGN EDFFHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.8900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0300 0.5100 1.4850 ;
        RECT  0.3600 1.0300 0.4800 1.5150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.7450 1.2550 11.0850 1.4650 ;
        RECT  10.7450 1.2300 11.0050 1.4650 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.0350 0.9900 11.4050 1.1100 ;
        RECT  10.5050 0.9700 11.2950 1.0900 ;
        RECT  11.0350 0.9400 11.2950 1.1100 ;
        RECT  10.7250 0.4100 10.8450 1.0900 ;
        RECT  10.0250 0.4100 10.8450 0.5300 ;
        RECT  10.0250 0.4100 10.1450 1.0100 ;
        RECT  10.0050 0.8900 10.1250 1.4600 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0450 0.8000 8.0450 0.9200 ;
        RECT  7.9250 0.6800 8.0450 0.9200 ;
        RECT  7.6250 1.4500 7.8650 1.5900 ;
        RECT  5.0450 1.4500 7.8650 1.5700 ;
        RECT  6.9650 0.6800 7.0850 0.9200 ;
        RECT  6.7850 1.4500 7.0250 1.5900 ;
        RECT  5.8850 1.4500 6.1250 1.5900 ;
        RECT  6.0050 0.6800 6.1250 0.9200 ;
        RECT  5.5800 1.1750 5.7300 1.5700 ;
        RECT  5.6100 0.8000 5.7300 1.5700 ;
        RECT  5.0450 1.4500 5.2850 1.5900 ;
        RECT  5.0450 0.6800 5.1650 0.9200 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.8900 0.1800 ;
        RECT  11.0650 -0.1800 11.1850 0.8200 ;
        RECT  9.3050 -0.1800 9.4250 0.6400 ;
        RECT  8.4050 0.4600 8.6450 0.5800 ;
        RECT  8.5250 -0.1800 8.6450 0.5800 ;
        RECT  7.3850 -0.1800 7.6250 0.3200 ;
        RECT  6.4250 -0.1800 6.6650 0.3200 ;
        RECT  5.4650 -0.1800 5.7050 0.3200 ;
        RECT  4.5650 -0.1800 4.6850 0.6800 ;
        RECT  2.7250 0.4300 2.9650 0.5500 ;
        RECT  2.8450 -0.1800 2.9650 0.5500 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.8900 2.7900 ;
        RECT  11.0050 1.8250 11.1250 2.7900 ;
        RECT  9.3050 2.1000 9.5450 2.2200 ;
        RECT  9.3050 2.1000 9.4250 2.7900 ;
        RECT  8.3450 2.1000 8.5850 2.2200 ;
        RECT  8.3450 2.1000 8.4650 2.7900 ;
        RECT  7.2050 1.9500 7.4450 2.0700 ;
        RECT  7.2050 1.9500 7.3250 2.7900 ;
        RECT  6.3050 1.9500 6.5450 2.0750 ;
        RECT  6.3050 1.9500 6.4250 2.7900 ;
        RECT  5.4650 1.9500 5.7050 2.0750 ;
        RECT  5.4650 1.9500 5.5850 2.7900 ;
        RECT  4.6250 1.9500 4.8650 2.0750 ;
        RECT  4.6250 1.9500 4.7450 2.7900 ;
        RECT  2.7250 1.7500 2.8450 2.7900 ;
        RECT  0.5550 1.6350 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6450 1.7050 11.6050 1.7050 11.6050 1.8250 11.4850 1.8250 11.4850 1.7050
                 10.5050 1.7050 10.5050 1.2400 10.6250 1.2400 10.6250 1.5850 11.5250 1.5850
                 11.5250 0.8200 11.4850 0.8200 11.4850 0.5800 11.6050 0.5800 11.6050 0.7000
                 11.6450 0.7000 ;
        POLYGON  10.6050 0.7700 10.4850 0.7700 10.4850 0.8500 10.3850 0.8500 10.3850 2.2100
                 10.2650 2.2100 10.2650 1.9800 8.2650 1.9800 8.2650 1.8300 4.4100 1.8300 4.4100 2.1700
                 4.1450 2.1700 4.1450 2.2300 2.9650 2.2300 2.9650 1.6300 2.5550 1.6300 2.5550 2.2300
                 1.5450 2.2300 1.5450 1.5900 1.4250 1.5900 1.4250 0.7200 1.3050 0.7200 1.3050 0.6000
                 1.5450 0.6000 1.5450 1.4700 1.6650 1.4700 1.6650 2.1100 2.4350 2.1100 2.4350 1.5100
                 3.0850 1.5100 3.0850 2.1100 4.0250 2.1100 4.0250 2.0500 4.2900 2.0500 4.2900 1.7100
                 8.3850 1.7100 8.3850 1.8600 10.2650 1.8600 10.2650 0.7300 10.3650 0.7300
                 10.3650 0.6500 10.6050 0.6500 ;
        POLYGON  10.0250 1.7400 9.7650 1.7400 9.7650 1.6200 9.0650 1.6200 9.0650 1.7400 8.8250 1.7400
                 8.8250 1.6200 8.8850 1.6200 8.8850 1.3300 7.0650 1.3300 7.0650 1.1300 7.3050 1.1300
                 7.3050 1.2100 8.8850 1.2100 8.8850 0.5900 9.0050 0.5900 9.0050 0.7600 9.6650 0.7600
                 9.6650 0.6500 9.9050 0.6500 9.9050 0.7700 9.7850 0.7700 9.7850 0.8800 9.0050 0.8800
                 9.0050 1.5000 9.8850 1.5000 9.8850 1.6200 10.0250 1.6200 ;
        POLYGON  8.7650 1.0900 8.5250 1.0900 8.5250 0.8200 8.1650 0.8200 8.1650 0.5600 4.9250 0.5600
                 4.9250 0.9200 4.4850 0.9200 4.4850 1.5900 4.1700 1.5900 4.1700 1.6500 4.1650 1.6500
                 4.1650 1.9300 3.9250 1.9300 3.9250 1.5300 4.0500 1.5300 4.0500 1.4700 4.3650 1.4700
                 4.3650 0.9200 3.9250 0.9200 3.9250 0.5400 4.0450 0.5400 4.0450 0.8000 4.8050 0.8000
                 4.8050 0.4400 8.2850 0.4400 8.2850 0.7000 8.6450 0.7000 8.6450 0.9700 8.7650 0.9700 ;
        POLYGON  4.2450 1.3500 4.1250 1.3500 4.1250 1.1600 3.6850 1.1600 3.6850 1.1200 3.5650 1.1200
                 3.5650 0.8800 3.6850 0.8800 3.6850 0.4800 3.2050 0.4800 3.2050 0.7900 2.3850 0.7900
                 2.3850 1.1200 2.2450 1.1200 2.2450 0.8800 2.2650 0.8800 2.2650 0.4800 1.7850 0.4800
                 1.7850 0.8400 1.8050 0.8400 1.8050 1.3500 1.6850 1.3500 1.6850 0.9600 1.6650 0.9600
                 1.6650 0.4800 1.1350 0.4800 1.1350 1.6350 1.0950 1.6350 1.0950 1.7550 0.9750 1.7550
                 0.9750 1.5150 1.0150 1.5150 1.0150 0.6700 0.9750 0.6700 0.9750 0.3600 2.6050 0.3600
                 2.6050 0.6700 3.0850 0.6700 3.0850 0.3600 3.8050 0.3600 3.8050 1.0400 4.2450 1.0400 ;
        POLYGON  3.5650 0.7200 3.4450 0.7200 3.4450 1.9900 3.3250 1.9900 3.3250 1.3900 2.7450 1.3900
                 2.7450 1.1500 2.8650 1.1500 2.8650 1.2700 3.3250 1.2700 3.3250 0.6000 3.5650 0.6000 ;
        POLYGON  3.2050 1.1500 3.0850 1.1500 3.0850 1.0300 2.6250 1.0300 2.6250 1.3600 2.1250 1.3600
                 2.1250 1.9900 2.0050 1.9900 2.0050 0.7200 1.9050 0.7200 1.9050 0.6000 2.1450 0.6000
                 2.1450 0.7200 2.1250 0.7200 2.1250 1.2400 2.5050 1.2400 2.5050 0.9100 3.2050 0.9100 ;
        POLYGON  0.8950 0.9500 0.6550 0.9500 0.6550 0.9100 0.2400 0.9100 0.2400 1.6350 0.2550 1.6350
                 0.2550 1.8750 0.1350 1.8750 0.1350 1.7550 0.1200 1.7550 0.1200 0.6700 0.1350 0.6700
                 0.1350 0.4300 0.2550 0.4300 0.2550 0.7900 0.8950 0.7900 ;
    END
END EDFFHQX8

MACRO EDFFHQX4
    CLASS CORE ;
    FOREIGN EDFFHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.1500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0600 0.5100 1.5150 ;
        RECT  0.3600 1.0300 0.4800 1.5150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0600 1.0300 9.2400 1.4500 ;
        RECT  9.1200 1.0100 9.2400 1.4500 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5850 1.2300 9.8450 1.3800 ;
        RECT  9.5000 1.1400 9.7050 1.2600 ;
        RECT  9.5000 0.7700 9.6200 1.2600 ;
        RECT  8.8200 0.7700 9.6200 0.8900 ;
        RECT  8.7000 0.9800 8.9400 1.1000 ;
        RECT  8.8200 0.3600 8.9400 1.1000 ;
        RECT  8.2200 0.3600 8.9400 0.4800 ;
        RECT  8.2200 0.3600 8.3400 1.0800 ;
        RECT  8.1800 0.9600 8.3000 1.4400 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.7944  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1450 0.6500 6.3850 0.7700 ;
        RECT  6.0250 1.5800 6.2650 1.7100 ;
        RECT  5.0650 0.9400 6.2650 1.0600 ;
        RECT  6.1450 0.6500 6.2650 1.0600 ;
        RECT  5.0650 1.5800 6.2650 1.7000 ;
        RECT  5.1250 1.4700 5.2450 1.7100 ;
        RECT  5.0650 0.6500 5.1850 1.7000 ;
        RECT  4.9450 1.5200 5.2450 1.6700 ;
        RECT  4.9450 0.6500 5.1850 0.7700 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.1500 0.1800 ;
        RECT  9.2600 -0.1800 9.3800 0.6500 ;
        RECT  7.6450 -0.1800 7.7650 0.4500 ;
        RECT  6.7450 -0.1800 6.8650 0.6400 ;
        RECT  5.5450 0.4600 5.7850 0.5800 ;
        RECT  5.6650 -0.1800 5.7850 0.5800 ;
        RECT  4.4650 -0.1800 4.5850 0.6800 ;
        RECT  2.6250 0.4300 2.8650 0.5500 ;
        RECT  2.7450 -0.1800 2.8650 0.5500 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.1500 2.7900 ;
        RECT  9.2600 1.8100 9.3800 2.7900 ;
        RECT  7.5250 2.1600 7.6450 2.7900 ;
        RECT  6.5650 2.0700 6.6850 2.7900 ;
        RECT  5.5450 2.0700 5.7850 2.1900 ;
        RECT  5.5450 2.0700 5.6650 2.7900 ;
        RECT  4.5850 2.0700 4.8250 2.1900 ;
        RECT  4.5850 2.0700 4.7050 2.7900 ;
        RECT  2.7450 1.7500 2.8650 2.7900 ;
        RECT  0.6150 2.1550 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.0850 1.6900 9.8600 1.6900 9.8600 1.8100 9.7400 1.8100 9.7400 1.6900 8.8200 1.6900
                 8.8200 1.4200 8.7000 1.4200 8.7000 1.3000 8.9400 1.3000 8.9400 1.5700 9.9650 1.5700
                 9.9650 1.0200 9.7400 1.0200 9.7400 0.6000 9.8600 0.6000 9.8600 0.9000 10.0850 0.9000 ;
        POLYGON  8.7000 0.8600 8.5800 0.8600 8.5800 2.2100 8.4600 2.2100 8.4600 2.0400 7.6650 2.0400
                 7.6650 1.9500 4.2150 1.9500 4.2150 2.2300 3.0350 2.2300 3.0350 1.6300 2.6250 1.6300
                 2.6250 2.2300 1.4450 2.2300 1.4450 1.5900 1.3450 1.5900 1.3450 0.7200 1.3050 0.7200
                 1.3050 0.6000 1.5450 0.6000 1.5450 0.7200 1.4650 0.7200 1.4650 1.4700 1.5650 1.4700
                 1.5650 2.1100 2.5050 2.1100 2.5050 1.5100 3.1550 1.5100 3.1550 2.1100 4.0950 2.1100
                 4.0950 1.8300 7.7850 1.8300 7.7850 1.9200 8.4600 1.9200 8.4600 0.7400 8.5800 0.7400
                 8.5800 0.6000 8.7000 0.6000 ;
        POLYGON  8.1600 1.8000 8.0400 1.8000 8.0400 1.6800 7.9400 1.6800 7.9400 1.5600 7.1650 1.5600
                 7.1650 1.7100 7.0450 1.7100 7.0450 1.4600 5.8850 1.4600 5.8850 1.2100 6.1250 1.2100
                 6.1250 1.3400 7.4050 1.3400 7.4050 0.7800 7.1650 0.7800 7.1650 0.5000 7.2850 0.5000
                 7.2850 0.6600 7.5250 0.6600 7.5250 0.7200 7.9800 0.7200 7.9800 0.6000 8.1000 0.6000
                 8.1000 0.8400 7.5250 0.8400 7.5250 1.4400 8.0600 1.4400 8.0600 1.5600 8.1600 1.5600 ;
        POLYGON  7.2850 1.0200 6.9450 1.0200 6.9450 1.2200 6.7050 1.2200 6.7050 1.1000 6.8250 1.1000
                 6.8250 0.8800 6.5050 0.8800 6.5050 0.5300 6.0250 0.5300 6.0250 0.8200 5.3050 0.8200
                 5.3050 0.5300 4.8250 0.5300 4.8250 0.9200 4.4650 0.9200 4.4650 1.6100 4.1250 1.6100
                 4.1250 1.7100 3.8850 1.7100 3.8850 1.5300 4.0050 1.5300 4.0050 1.4900 4.3450 1.4900
                 4.3450 0.9200 3.8250 0.9200 3.8250 0.5400 3.9450 0.5400 3.9450 0.8000 4.7050 0.8000
                 4.7050 0.4100 5.4250 0.4100 5.4250 0.7000 5.9050 0.7000 5.9050 0.4100 6.6250 0.4100
                 6.6250 0.7600 6.9450 0.7600 6.9450 0.9000 7.2850 0.9000 ;
        POLYGON  4.2250 1.3700 4.1050 1.3700 4.1050 1.2500 3.5850 1.2500 3.5850 1.1200 3.5650 1.1200
                 3.5650 0.8800 3.5850 0.8800 3.5850 0.4800 3.1050 0.4800 3.1050 0.7900 2.3850 0.7900
                 2.3850 1.1200 2.1450 1.1200 2.1450 0.8800 2.2650 0.8800 2.2650 0.4800 1.7850 0.4800
                 1.7850 0.9600 1.7050 0.9600 1.7050 1.3500 1.5850 1.3500 1.5850 0.8400 1.6650 0.8400
                 1.6650 0.4800 1.1850 0.4800 1.1850 1.6350 1.1750 1.6350 1.1750 1.7550 1.0550 1.7550
                 1.0550 1.5150 1.0650 1.5150 1.0650 0.6700 0.9750 0.6700 0.9750 0.3600 2.5050 0.3600
                 2.5050 0.6700 2.9850 0.6700 2.9850 0.3600 3.7050 0.3600 3.7050 1.1300 4.2250 1.1300 ;
        POLYGON  3.4650 0.7200 3.4450 0.7200 3.4450 1.3900 3.3950 1.3900 3.3950 1.9900 3.2750 1.9900
                 3.2750 1.3900 2.7450 1.3900 2.7450 1.1500 2.8650 1.1500 2.8650 1.2700 3.3250 1.2700
                 3.3250 0.7200 3.2250 0.7200 3.2250 0.6000 3.4650 0.6000 ;
        POLYGON  3.2050 1.1500 3.0850 1.1500 3.0850 1.0300 2.6250 1.0300 2.6250 1.3600 2.0250 1.3600
                 2.0250 1.9900 1.9050 1.9900 1.9050 0.6000 2.1450 0.6000 2.1450 0.7200 2.0250 0.7200
                 2.0250 1.2400 2.5050 1.2400 2.5050 0.9100 3.2050 0.9100 ;
        POLYGON  0.9450 0.9500 0.7050 0.9500 0.7050 0.9100 0.2400 0.9100 0.2400 1.6350 0.2550 1.6350
                 0.2550 1.8750 0.1350 1.8750 0.1350 1.7550 0.1200 1.7550 0.1200 0.6700 0.1350 0.6700
                 0.1350 0.4300 0.2550 0.4300 0.2550 0.7900 0.9450 0.7900 ;
    END
END EDFFHQX4

MACRO EDFFHQX2
    CLASS CORE ;
    FOREIGN EDFFHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.2300 0.8550 1.4000 ;
        RECT  0.4700 1.2300 0.8550 1.3850 ;
        RECT  0.4700 1.1100 0.5900 1.3850 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8200 1.1300 8.0600 1.3350 ;
        RECT  7.9000 1.0800 8.0500 1.4750 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1900 0.8400 8.3400 1.1450 ;
        RECT  7.1600 0.8400 8.3400 0.9600 ;
        RECT  7.3200 0.3600 7.4400 0.9600 ;
        RECT  6.6800 0.3600 7.4400 0.4800 ;
        RECT  7.1600 0.8400 7.2800 1.1700 ;
        RECT  6.6800 0.3600 6.8000 1.2700 ;
        RECT  6.5800 1.1500 6.7000 1.3900 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.4200 1.5300 5.6600 1.6500 ;
        RECT  5.4200 0.6700 5.6600 0.7900 ;
        RECT  5.4200 0.6700 5.5400 1.6500 ;
        RECT  5.2900 1.1750 5.5400 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.6600 -0.1800 7.7800 0.6600 ;
        RECT  6.0200 -0.1800 6.1400 0.6600 ;
        RECT  4.9400 -0.1800 5.0600 0.6800 ;
        RECT  2.9600 0.4900 3.2000 0.6100 ;
        RECT  2.9600 -0.1800 3.0800 0.6100 ;
        RECT  0.5900 0.5700 0.8300 0.6900 ;
        RECT  0.5900 -0.1800 0.7100 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  8.0200 1.8350 8.1400 2.7900 ;
        RECT  5.9000 2.0100 6.1400 2.1300 ;
        RECT  5.9000 2.0100 6.0200 2.7900 ;
        RECT  4.9400 2.0100 5.1800 2.1300 ;
        RECT  4.9400 2.0100 5.0600 2.7900 ;
        RECT  3.0200 1.7200 3.1400 2.7900 ;
        RECT  2.9000 1.7200 3.1400 1.9300 ;
        RECT  0.6500 1.5700 0.7700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.5800 1.8350 8.5600 1.8350 8.5600 2.0000 8.4400 2.0000 8.4400 1.7150 7.5200 1.7150
                 7.5200 1.1500 7.6400 1.1500 7.6400 1.5950 8.4600 1.5950 8.4600 0.7200 8.3800 0.7200
                 8.3800 0.4800 8.5000 0.4800 8.5000 0.6000 8.5800 0.6000 ;
        POLYGON  7.2000 0.7200 7.0400 0.7200 7.0400 2.1200 6.9200 2.1200 6.9200 1.8900 4.7050 1.8900
                 4.7050 2.2300 3.2600 2.2300 3.2600 1.6000 2.7800 1.6000 2.7800 2.2300 1.6600 2.2300
                 1.6600 1.5900 1.5000 1.5900 1.5000 0.7200 1.4000 0.7200 1.4000 0.6000 1.6400 0.6000
                 1.6400 0.7200 1.6200 0.7200 1.6200 1.4700 1.7800 1.4700 1.7800 2.1100 2.6600 2.1100
                 2.6600 1.4800 3.3800 1.4800 3.3800 2.1100 4.5850 2.1100 4.5850 1.7700 6.9200 1.7700
                 6.9200 0.6000 7.2000 0.6000 ;
        POLYGON  6.6200 1.6500 6.3400 1.6500 6.3400 1.4100 5.7400 1.4100 5.7400 1.1500 5.8600 1.1500
                 5.8600 1.2900 6.3400 1.2900 6.3400 0.7300 6.4400 0.7300 6.4400 0.6100 6.5600 0.6100
                 6.5600 0.8500 6.4600 0.8500 6.4600 1.5300 6.6200 1.5300 ;
        POLYGON  6.2200 1.1700 6.1000 1.1700 6.1000 0.9000 5.7800 0.9000 5.7800 0.5500 5.3000 0.5500
                 5.3000 0.9200 4.8000 0.9200 4.8000 1.6300 4.3200 1.6300 4.3200 1.9900 4.2000 1.9900
                 4.2000 1.4700 4.3200 1.4700 4.3200 1.5100 4.6800 1.5100 4.6800 0.9200 4.1600 0.9200
                 4.1600 0.5400 4.2800 0.5400 4.2800 0.8000 5.1800 0.8000 5.1800 0.4300 5.9000 0.4300
                 5.9000 0.7800 6.2200 0.7800 ;
        POLYGON  4.5600 1.3900 4.4400 1.3900 4.4400 1.1600 3.9200 1.1600 3.9200 1.0400 3.8000 1.0400
                 3.8000 0.9200 3.9200 0.9200 3.9200 0.4800 3.4400 0.4800 3.4400 0.8500 2.6250 0.8500
                 2.6250 0.4800 2.4800 0.4800 2.4800 1.1200 2.3600 1.1200 2.3600 0.4800 1.8800 0.4800
                 1.8800 1.2100 1.9800 1.2100 1.9800 1.3300 1.7400 1.3300 1.7400 1.2100 1.7600 1.2100
                 1.7600 0.4800 1.1900 0.4800 1.1900 0.6300 1.2300 0.6300 1.2300 1.5700 1.1900 1.5700
                 1.1900 1.6900 1.0700 1.6900 1.0700 1.4500 1.1100 1.4500 1.1100 0.7500 1.0700 0.7500
                 1.0700 0.3600 2.7450 0.3600 2.7450 0.7300 3.3200 0.7300 3.3200 0.3600 4.0400 0.3600
                 4.0400 1.0400 4.5600 1.0400 ;
        POLYGON  3.8000 0.7200 3.6800 0.7200 3.6800 1.3300 3.6200 1.3300 3.6200 1.9900 3.5000 1.9900
                 3.5000 1.3300 2.8400 1.3300 2.8400 1.2100 3.5600 1.2100 3.5600 0.6000 3.8000 0.6000 ;
        POLYGON  3.4400 1.0900 2.7200 1.0900 2.7200 1.3600 2.2400 1.3600 2.2400 1.9900 2.1200 1.9900
                 2.1200 0.7200 2.0000 0.7200 2.0000 0.6000 2.2400 0.6000 2.2400 1.2400 2.6000 1.2400
                 2.6000 0.9700 3.4400 0.9700 ;
        POLYGON  0.9900 1.0100 0.7500 1.0100 0.7500 0.9900 0.3500 0.9900 0.3500 1.6900 0.2300 1.6900
                 0.2300 0.5100 0.3500 0.5100 0.3500 0.8700 0.9900 0.8700 ;
    END
END EDFFHQX2

MACRO EDFFHQX1
    CLASS CORE ;
    FOREIGN EDFFHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0900 0.5100 1.5450 ;
        RECT  0.3600 1.0700 0.4800 1.5450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.2300 7.5250 1.4600 ;
        RECT  7.2750 1.0800 7.3950 1.4900 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5550 0.9400 7.8150 1.0900 ;
        RECT  7.5550 0.9400 7.7950 1.1100 ;
        RECT  6.9450 0.8400 7.6750 0.9600 ;
        RECT  7.1050 0.3600 7.2250 0.9600 ;
        RECT  6.3450 0.3600 7.2250 0.4800 ;
        RECT  6.9450 0.8400 7.0650 1.1500 ;
        RECT  6.3450 0.3600 6.4650 1.4600 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0850 1.5300 5.4050 1.6500 ;
        RECT  5.0850 0.6300 5.2050 1.6500 ;
        RECT  5.0000 1.1750 5.2050 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.4450 -0.1800 7.5650 0.7200 ;
        RECT  5.5650 -0.1800 5.6850 0.7300 ;
        RECT  4.4850 0.5000 4.7250 0.6200 ;
        RECT  4.4850 -0.1800 4.6050 0.6200 ;
        RECT  2.7050 0.4300 2.9450 0.5500 ;
        RECT  2.7050 -0.1800 2.8250 0.5500 ;
        RECT  0.5550 -0.1800 0.6750 0.7100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.3850 1.8500 7.5050 2.7900 ;
        RECT  5.6250 2.1000 5.8650 2.2200 ;
        RECT  5.6250 2.1000 5.7450 2.7900 ;
        RECT  4.6850 2.0100 4.9250 2.1300 ;
        RECT  4.6850 2.0100 4.8050 2.7900 ;
        RECT  2.7950 1.7500 2.9150 2.7900 ;
        RECT  0.5550 1.6650 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.0550 1.7300 7.9850 1.7300 7.9850 1.8500 7.8650 1.8500 7.8650 1.7300 6.9450 1.7300
                 6.9450 1.4200 6.8250 1.4200 6.8250 1.3000 7.0650 1.3000 7.0650 1.6100 7.9350 1.6100
                 7.9350 0.7200 7.8650 0.7200 7.8650 0.4800 7.9850 0.4800 7.9850 0.6000 8.0550 0.6000 ;
        POLYGON  6.9850 0.7200 6.7050 0.7200 6.7050 1.5600 6.7650 1.5600 6.7650 2.2100 6.6450 2.2100
                 6.6450 1.9800 5.8500 1.9800 5.8500 1.8900 4.3800 1.8900 4.3800 2.2300 3.0850 2.2300
                 3.0850 1.6300 2.6750 1.6300 2.6750 2.2300 1.5250 2.2300 1.5250 1.5900 1.3650 1.5900
                 1.3650 0.7200 1.3050 0.7200 1.3050 0.6000 1.5450 0.6000 1.5450 0.7200 1.4850 0.7200
                 1.4850 1.4700 1.6450 1.4700 1.6450 2.1100 2.5550 2.1100 2.5550 1.5100 3.2050 1.5100
                 3.2050 2.1100 4.2600 2.1100 4.2600 1.7700 5.9700 1.7700 5.9700 1.8600 6.6450 1.8600
                 6.6450 1.6800 6.5850 1.6800 6.5850 0.6000 6.9850 0.6000 ;
        POLYGON  6.4050 1.7400 6.0900 1.7400 6.0900 1.4100 5.5050 1.4100 5.5050 1.2900 6.0900 1.2900
                 6.0900 0.7700 5.9850 0.7700 5.9850 0.6500 6.2250 0.6500 6.2250 0.7700 6.2100 0.7700
                 6.2100 1.6200 6.4050 1.6200 ;
        POLYGON  5.9650 1.0900 5.7250 1.0900 5.7250 0.9700 5.3250 0.9700 5.3250 0.5100 4.9650 0.5100
                 4.9650 0.8600 4.5450 0.8600 4.5450 1.6300 4.0650 1.6300 4.0650 1.9900 3.9450 1.9900
                 3.9450 1.4700 4.0650 1.4700 4.0650 1.5100 4.4250 1.5100 4.4250 0.8600 3.9250 0.8600
                 3.9250 0.7800 3.9050 0.7800 3.9050 0.5400 4.0250 0.5400 4.0250 0.6600 4.0450 0.6600
                 4.0450 0.7400 4.8450 0.7400 4.8450 0.3900 5.4450 0.3900 5.4450 0.8500 5.8450 0.8500
                 5.8450 0.9700 5.9650 0.9700 ;
        POLYGON  4.3050 1.3900 4.1850 1.3900 4.1850 1.1000 3.6650 1.1000 3.6650 1.0600 3.5650 1.0600
                 3.5650 0.9400 3.6650 0.9400 3.6650 0.4800 3.1850 0.4800 3.1850 0.7900 2.3850 0.7900
                 2.3850 1.1200 2.2250 1.1200 2.2250 0.8800 2.2650 0.8800 2.2650 0.4800 1.7850 0.4800
                 1.7850 1.2100 1.8450 1.2100 1.8450 1.3300 1.6050 1.3300 1.6050 1.2100 1.6650 1.2100
                 1.6650 0.4800 1.1350 0.4800 1.1350 1.6650 1.0950 1.6650 1.0950 1.7850 0.9750 1.7850
                 0.9750 1.5450 1.0150 1.5450 1.0150 0.7100 0.9750 0.7100 0.9750 0.3600 2.5850 0.3600
                 2.5850 0.6700 3.0650 0.6700 3.0650 0.3600 3.7850 0.3600 3.7850 0.9400 3.8050 0.9400
                 3.8050 0.9800 4.3050 0.9800 ;
        POLYGON  3.5450 0.7200 3.4450 0.7200 3.4450 1.9900 3.3250 1.9900 3.3250 1.3900 2.7450 1.3900
                 2.7450 1.1500 2.8650 1.1500 2.8650 1.2700 3.3250 1.2700 3.3250 0.7200 3.3050 0.7200
                 3.3050 0.6000 3.5450 0.6000 ;
        POLYGON  3.2050 1.1500 3.0850 1.1500 3.0850 1.0300 2.6250 1.0300 2.6250 1.3600 2.1050 1.3600
                 2.1050 1.9900 1.9850 1.9900 1.9850 0.7200 1.9050 0.7200 1.9050 0.6000 2.1450 0.6000
                 2.1450 0.7200 2.1050 0.7200 2.1050 1.2400 2.5050 1.2400 2.5050 0.9100 3.2050 0.9100 ;
        POLYGON  0.8950 0.9900 0.6550 0.9900 0.6550 0.9500 0.2400 0.9500 0.2400 1.6650 0.2550 1.6650
                 0.2550 1.9050 0.1350 1.9050 0.1350 1.7850 0.1200 1.7850 0.1200 0.7100 0.1350 0.7100
                 0.1350 0.4700 0.2550 0.4700 0.2550 0.8300 0.8950 0.8300 ;
    END
END EDFFHQX1

MACRO DLY4X4
    CLASS CORE ;
    FOREIGN DLY4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9950 1.4000 2.2350 1.5200 ;
        RECT  2.0550 0.5900 2.1750 1.5200 ;
        RECT  1.2300 1.0250 2.1750 1.1450 ;
        RECT  1.2150 0.8850 1.3800 1.0250 ;
        RECT  1.0350 1.4000 1.3500 1.5200 ;
        RECT  1.2300 0.8850 1.3500 1.5200 ;
        RECT  1.2150 0.5900 1.3350 1.0250 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.2500 10.5750 1.4900 ;
        RECT  10.2500 1.3700 10.5750 1.4900 ;
        RECT  10.2200 1.4650 10.3700 1.7250 ;
        END
    END A
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.2350 -0.1800 10.3550 0.8900 ;
        RECT  9.6850 1.2400 9.9550 1.3600 ;
        RECT  9.8350 -0.1800 9.9550 1.3600 ;
        RECT  9.6850 1.2400 9.8050 1.4800 ;
        RECT  8.3650 -0.1800 8.4850 0.3800 ;
        RECT  7.5850 -0.1800 7.7050 1.3600 ;
        RECT  7.4850 1.2400 7.6050 1.4800 ;
        RECT  6.6350 1.2000 6.8750 1.3200 ;
        RECT  6.7150 -0.1800 6.8350 1.3200 ;
        RECT  6.0150 -0.1800 6.1350 0.8400 ;
        RECT  5.1550 1.5100 5.4150 1.6300 ;
        RECT  5.1550 -0.1800 5.2750 1.6300 ;
        RECT  4.1350 1.4800 4.5550 1.7200 ;
        RECT  4.4350 0.9800 4.5550 1.7200 ;
        RECT  4.2250 0.9800 4.5550 1.1000 ;
        RECT  4.2250 -0.1800 4.3450 1.1000 ;
        RECT  3.8850 -0.1800 4.0050 0.8600 ;
        RECT  3.0750 1.0000 3.1950 1.2400 ;
        RECT  2.8150 1.0000 3.1950 1.1200 ;
        RECT  2.8150 -0.1800 2.9350 1.1200 ;
        RECT  2.4750 -0.1800 2.5950 0.6400 ;
        RECT  1.6350 -0.1800 1.7550 0.6400 ;
        RECT  0.7950 -0.1800 0.9150 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.2450 2.2300 10.3650 2.7900 ;
        RECT  8.9450 1.0000 9.0650 1.2400 ;
        RECT  7.8250 1.0000 9.0650 1.1200 ;
        RECT  8.4250 1.6800 8.5450 2.7900 ;
        RECT  7.9650 1.0000 8.0850 2.7900 ;
        RECT  7.8250 1.0000 8.0850 1.2400 ;
        RECT  6.1950 2.1600 6.3150 2.7900 ;
        RECT  6.0750 2.1600 6.3150 2.2800 ;
        RECT  4.9950 1.7900 5.1150 2.7900 ;
        RECT  3.5150 2.0800 3.7550 2.2000 ;
        RECT  3.5150 2.0800 3.6350 2.7900 ;
        RECT  2.5350 1.8800 2.6550 2.7900 ;
        RECT  1.5150 1.8800 1.7550 2.0000 ;
        RECT  1.5150 1.8800 1.6350 2.7900 ;
        RECT  0.5550 1.8800 0.7950 2.0000 ;
        RECT  0.5550 1.8800 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.8450 1.8500 10.7250 1.8500 10.7250 1.7300 10.6950 1.7300 10.6950 1.1300
                 10.3350 1.1300 10.3350 1.1700 10.0750 1.1700 10.0750 1.0500 10.2150 1.0500
                 10.2150 1.0100 10.6550 1.0100 10.6550 0.6500 10.7750 0.6500 10.7750 0.8900
                 10.8150 0.8900 10.8150 1.6100 10.8450 1.6100 ;
        POLYGON  9.7150 0.8900 9.5650 0.8900 9.5650 1.6000 9.6650 1.6000 9.6650 1.8400 9.5450 1.8400
                 9.5450 1.7200 9.4450 1.7200 9.4450 0.7700 9.5950 0.7700 9.5950 0.6500 9.5600 0.6500
                 9.5600 0.5400 8.7650 0.5400 8.7650 0.5200 8.6450 0.5200 8.6450 0.4000 8.8850 0.4000
                 8.8850 0.4200 9.6800 0.4200 9.6800 0.5300 9.7150 0.5300 ;
        POLYGON  9.3250 1.4800 9.1850 1.4800 9.1850 1.8000 9.0650 1.8000 9.0650 1.4800 8.2050 1.4800
                 8.2050 1.2400 8.3250 1.2400 8.3250 1.3600 9.2050 1.3600 9.2050 0.6600 9.3250 0.6600 ;
        POLYGON  7.8450 1.8000 6.0550 1.8000 6.0550 1.7700 6.0150 1.7700 6.0150 1.5300 6.0550 1.5300
                 6.0550 0.9600 6.2950 0.9600 6.2950 0.3600 6.5350 0.3600 6.5350 1.0800 6.1750 1.0800
                 6.1750 1.6800 7.2450 1.6800 7.2450 0.7800 7.3450 0.7800 7.3450 0.6600 7.4650 0.6600
                 7.4650 0.9000 7.3650 0.9000 7.3650 1.6800 7.8450 1.6800 ;
        POLYGON  7.1150 1.5600 6.2950 1.5600 6.2950 1.4400 6.9950 1.4400 6.9950 1.0800 6.9550 1.0800
                 6.9550 0.6200 7.0750 0.6200 7.0750 0.9600 7.1150 0.9600 ;
        POLYGON  7.0150 2.0400 5.7750 2.0400 5.7750 0.4800 5.3950 0.4800 5.3950 0.3600 5.8950 0.3600
                 5.8950 1.9200 7.0150 1.9200 ;
        POLYGON  5.6550 1.8700 5.5550 1.8700 5.5550 2.0900 5.4350 2.0900 5.4350 1.7500 5.5350 1.7500
                 5.5350 1.1300 5.6550 1.1300 ;
        POLYGON  5.0350 0.8600 4.9150 0.8600 4.9150 0.4800 4.7750 0.4800 4.7750 0.3600 5.0350 0.3600 ;
        POLYGON  4.7950 1.9700 4.3950 1.9700 4.3950 2.0900 4.2750 2.0900 4.2750 1.9700 4.2600 1.9700
                 4.2600 1.9600 2.8150 1.9600 2.8150 1.8400 4.3800 1.8400 4.3800 1.8500 4.6750 1.8500
                 4.6750 0.8000 4.4650 0.8000 4.4650 0.6800 4.7950 0.6800 ;
        POLYGON  4.3150 1.3400 3.5550 1.3400 3.5550 0.9400 3.6750 0.9400 3.6750 1.2200 4.3150 1.2200 ;
        POLYGON  3.4950 1.7200 2.6950 1.7200 2.6950 1.7600 0.6150 1.7600 0.6150 1.0000 0.7350 1.0000
                 0.7350 1.6400 2.5750 1.6400 2.5750 1.6000 3.3150 1.6000 3.3150 0.8800 3.1750 0.8800
                 3.1750 0.5800 3.0550 0.5800 3.0550 0.4600 3.2950 0.4600 3.2950 0.7600 3.4350 0.7600
                 3.4350 1.4600 3.4950 1.4600 ;
        POLYGON  1.0750 1.1700 0.9550 1.1700 0.9550 0.8800 0.4950 0.8800 0.4950 1.4600 0.2550 1.4600
                 0.2550 1.9900 0.1350 1.9900 0.1350 1.3400 0.3750 1.3400 0.3750 0.5900 0.4950 0.5900
                 0.4950 0.7600 1.0750 0.7600 ;
    END
END DLY4X4

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.1500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.6400 1.1650 9.7900 1.6150 ;
        RECT  9.6400 1.1650 9.7600 1.6400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8750 0.9400 1.1450 1.0900 ;
        RECT  0.8750 0.6800 0.9950 1.9900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.1500 0.1800 ;
        RECT  9.4750 -0.1800 9.5950 0.7650 ;
        RECT  9.0750 -0.1800 9.1950 1.0050 ;
        RECT  8.9750 0.8850 9.0950 1.4800 ;
        RECT  7.6050 -0.1800 7.7250 0.3800 ;
        RECT  6.7150 1.3000 6.9550 1.4200 ;
        RECT  6.8350 -0.1800 6.9550 1.4200 ;
        RECT  5.8750 1.2400 6.1150 1.3600 ;
        RECT  5.9650 -0.1800 6.0850 1.3600 ;
        RECT  5.3250 -0.1800 5.4450 0.3800 ;
        RECT  4.5850 -0.1800 4.7050 1.0900 ;
        RECT  4.5550 0.9700 4.6750 1.7700 ;
        RECT  3.6550 1.5900 3.9350 1.7100 ;
        RECT  3.6550 -0.1800 3.7750 1.7100 ;
        RECT  3.1950 -0.1800 3.3150 0.5300 ;
        RECT  2.7250 1.2000 2.8450 1.4400 ;
        RECT  2.6850 -0.1800 2.8050 1.3200 ;
        RECT  1.8850 -0.1800 2.0050 0.9200 ;
        RECT  0.3950 -0.1800 0.5150 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.1500 2.7900 ;
        RECT  9.4750 1.7600 9.5950 2.7900 ;
        RECT  8.2050 1.0000 8.3250 1.2400 ;
        RECT  7.0750 1.0400 8.3250 1.1600 ;
        RECT  7.6950 2.2000 7.8150 2.7900 ;
        RECT  7.2950 1.0400 7.4150 2.7900 ;
        RECT  5.3150 2.2000 5.5550 2.7900 ;
        RECT  4.2950 1.0400 4.4150 2.7900 ;
        RECT  4.1750 1.0400 4.4150 1.1600 ;
        RECT  3.1350 2.0800 3.3750 2.2000 ;
        RECT  3.2350 2.0800 3.3550 2.7900 ;
        RECT  2.3250 1.0400 2.5650 1.1800 ;
        RECT  1.5050 1.0400 2.5650 1.1600 ;
        RECT  1.5050 2.2800 1.9250 2.7900 ;
        RECT  1.5050 1.0400 1.6250 2.7900 ;
        RECT  0.4550 1.3400 0.5750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.0300 1.8800 10.0150 1.8800 10.0150 2.0000 9.8950 2.0000 9.8950 1.7600 9.9100 1.7600
                 9.9100 1.0450 9.3150 1.0450 9.3150 0.9250 9.8950 0.9250 9.8950 0.5250 10.0150 0.5250
                 10.0150 0.8050 10.0300 0.8050 ;
        POLYGON  8.9550 0.7650 8.8550 0.7650 8.8550 1.6400 8.9550 1.6400 8.9550 1.8800 8.8350 1.8800
                 8.8350 1.7600 8.7350 1.7600 8.7350 0.6450 8.8350 0.6450 8.8350 0.5250 8.8000 0.5250
                 8.8000 0.5200 7.8850 0.5200 7.8850 0.4000 8.9200 0.4000 8.9200 0.4050 8.9550 0.4050 ;
        POLYGON  8.5650 1.4800 8.4850 1.4800 8.4850 1.8000 8.3650 1.8000 8.3650 1.4800 7.5350 1.4800
                 7.5350 1.3000 7.7750 1.3000 7.7750 1.3600 8.4450 1.3600 8.4450 0.6600 8.5650 0.6600 ;
        POLYGON  7.1750 1.8400 5.2950 1.8400 5.2950 1.7500 5.2750 1.7500 5.2750 1.5100 5.2950 1.5100
                 5.2950 0.5000 5.6050 0.5000 5.6050 0.4000 5.8450 0.4000 5.8450 0.6200 5.4150 0.6200
                 5.4150 1.7200 6.4750 1.7200 6.4750 0.7800 6.5950 0.7800 6.5950 0.6600 6.7150 0.6600
                 6.7150 0.9000 6.5950 0.9000 6.5950 1.7200 7.1750 1.7200 ;
        POLYGON  6.3550 1.6000 5.5350 1.6000 5.5350 1.4800 6.2350 1.4800 6.2350 1.1200 6.2050 1.1200
                 6.2050 0.6600 6.3250 0.6600 6.3250 1.0000 6.3550 1.0000 ;
        POLYGON  6.2550 2.0800 5.0350 2.0800 5.0350 1.0900 4.9450 1.0900 4.9450 0.4800 4.8250 0.4800
                 4.8250 0.3600 5.0650 0.3600 5.0650 0.9700 5.1550 0.9700 5.1550 1.9600 6.2550 1.9600 ;
        POLYGON  4.9150 2.0100 4.7950 2.0100 4.7950 2.1300 4.6750 2.1300 4.6750 1.8900 4.7950 1.8900
                 4.7950 1.2100 4.9150 1.2100 ;
        POLYGON  4.4650 0.8400 4.2250 0.8400 4.2250 0.4800 4.1450 0.4800 4.1450 0.3600 4.3850 0.3600
                 4.3850 0.4800 4.3450 0.4800 4.3450 0.7200 4.4650 0.7200 ;
        POLYGON  4.1750 1.9700 4.0150 1.9700 4.0150 2.0900 3.8950 2.0900 3.8950 1.9700 3.7350 1.9700
                 3.7350 1.9600 2.7950 1.9600 2.7950 2.1600 2.0250 2.1600 2.0250 2.0400 2.6750 2.0400
                 2.6750 1.8400 3.8550 1.8400 3.8550 1.8500 4.0550 1.8500 4.0550 1.4700 3.9350 1.4700
                 3.9350 0.8600 3.8950 0.8600 3.8950 0.6200 4.0150 0.6200 4.0150 0.7400 4.0550 0.7400
                 4.0550 1.3500 4.1750 1.3500 ;
        POLYGON  3.0850 1.7200 2.5250 1.7200 2.5250 1.6800 2.4450 1.6800 2.4450 1.4200 1.7450 1.4200
                 1.7450 1.2800 1.9850 1.2800 1.9850 1.3000 2.5650 1.3000 2.5650 1.5600 2.9650 1.5600
                 2.9650 0.9200 2.9250 0.9200 2.9250 0.6800 3.0450 0.6800 3.0450 0.8000 3.0850 0.8000 ;
        POLYGON  1.5850 0.9200 1.3850 0.9200 1.3850 1.7800 1.2650 1.7800 1.2650 0.8000 1.4650 0.8000
                 1.4650 0.6800 1.4300 0.6800 1.4300 0.5600 0.7550 0.5600 0.7550 1.1800 0.5150 1.1800
                 0.5150 1.0600 0.6350 1.0600 0.6350 0.4400 1.5500 0.4400 1.5500 0.5600 1.5850 0.5600 ;
    END
END DLY4X1

MACRO DLY3X4
    CLASS CORE ;
    FOREIGN DLY3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3150 0.6800 5.5550 0.8000 ;
        RECT  5.3750 0.6800 5.4950 2.2100 ;
        RECT  4.4200 0.8850 5.4950 1.0050 ;
        RECT  5.3150 0.6800 5.4950 1.0050 ;
        RECT  4.5350 0.8850 4.6550 2.2100 ;
        RECT  4.4200 0.6800 4.5950 1.1450 ;
        RECT  4.3550 0.6800 4.5950 0.8000 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6600 0.8850 2.8600 1.1450 ;
        RECT  2.6050 1.0250 2.7800 1.2650 ;
        END
    END A
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.5700 0.9200 8.6900 1.7400 ;
        RECT  8.4350 0.9200 8.6900 1.0400 ;
        RECT  8.4350 -0.1800 8.5550 1.0400 ;
        RECT  7.7350 0.6000 7.9750 0.7200 ;
        RECT  7.8350 -0.1800 7.9550 0.7200 ;
        RECT  6.4550 1.2400 6.6350 1.4800 ;
        RECT  6.5150 -0.1800 6.6350 1.4800 ;
        RECT  5.9150 0.6800 6.1550 0.8000 ;
        RECT  5.9150 -0.1800 6.0350 0.8000 ;
        RECT  4.8350 -0.1800 5.0750 0.3200 ;
        RECT  3.8750 -0.1800 3.9950 0.5300 ;
        RECT  3.6250 1.0400 3.7450 1.4200 ;
        RECT  3.3150 1.0400 3.7450 1.1600 ;
        RECT  3.3150 -0.1800 3.4350 1.1600 ;
        RECT  2.5950 -0.1800 2.8350 0.3400 ;
        RECT  1.6550 1.3700 1.8950 1.4900 ;
        RECT  1.7750 0.7600 1.8950 1.4900 ;
        RECT  1.5750 0.7600 1.8950 0.8800 ;
        RECT  1.5750 -0.1800 1.6950 0.8800 ;
        RECT  1.1750 -0.1800 1.2950 0.6400 ;
        RECT  0.3750 -0.1800 0.4950 1.3600 ;
        RECT  0.3550 1.2400 0.4750 1.4800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.3300 1.1600 8.4500 1.4000 ;
        RECT  7.3700 1.1600 8.4500 1.2800 ;
        RECT  7.3700 1.7600 7.6100 2.7900 ;
        RECT  7.3700 1.0800 7.4900 2.7900 ;
        RECT  7.2350 1.0800 7.4900 1.2000 ;
        RECT  5.7950 1.5800 5.9150 2.7900 ;
        RECT  4.9550 1.5600 5.0750 2.7900 ;
        RECT  4.1150 1.9300 4.2350 2.7900 ;
        RECT  3.2250 1.2800 3.4650 1.4000 ;
        RECT  3.2250 1.2800 3.3450 2.7900 ;
        RECT  2.7850 1.6600 2.9050 2.7900 ;
        RECT  0.6150 1.0000 1.6550 1.1200 ;
        RECT  1.1750 1.6100 1.5350 1.7300 ;
        RECT  1.4150 1.0000 1.5350 1.7300 ;
        RECT  0.9750 1.8400 1.2950 2.7900 ;
        RECT  1.1750 1.6100 1.2950 2.7900 ;
        RECT  0.8550 1.8400 1.2950 1.9600 ;
        RECT  0.6150 0.7800 0.8550 1.1200 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.9300 2.0200 8.4100 2.0200 8.4100 1.9800 8.3300 1.9800 8.3300 1.6400 7.6900 1.6400
                 7.6900 1.4000 7.9300 1.4000 7.9300 1.5200 8.4500 1.5200 8.4500 1.8600 8.8100 1.8600
                 8.8100 0.8000 8.6750 0.8000 8.6750 0.6800 8.9300 0.6800 ;
        POLYGON  8.3150 0.4800 8.2150 0.4800 8.2150 0.9600 7.4950 0.9600 7.4950 0.6200 6.8750 0.6200
                 6.8750 1.7200 6.5550 1.7200 6.5550 1.8400 6.4350 1.8400 6.4350 1.6000 6.7550 1.6000
                 6.7550 0.5000 7.6150 0.5000 7.6150 0.8400 8.0950 0.8400 8.0950 0.4800 8.0750 0.4800
                 8.0750 0.3600 8.3150 0.3600 ;
        POLYGON  7.3750 0.8600 7.2550 0.8600 7.2550 0.9600 7.1150 0.9600 7.1150 1.5600 7.1900 1.5600
                 7.1900 2.2100 7.0700 2.2100 7.0700 2.0800 6.0350 2.0800 6.0350 1.4200 5.6150 1.4200
                 5.6150 1.3000 6.1550 1.3000 6.1550 1.9600 6.9950 1.9600 6.9950 0.8400 7.1350 0.8400
                 7.1350 0.7400 7.3750 0.7400 ;
        POLYGON  6.3950 1.0400 5.6750 1.0400 5.6750 0.5600 4.2350 0.5600 4.2350 0.7700 3.9850 0.7700
                 3.9850 1.6600 3.9050 1.6600 3.9050 1.7800 3.7850 1.7800 3.7850 1.5400 3.8650 1.5400
                 3.8650 0.9200 3.5550 0.9200 3.5550 0.6500 4.1150 0.6500 4.1150 0.4400 5.7950 0.4400
                 5.7950 0.9200 6.2750 0.9200 6.2750 0.4800 6.1550 0.4800 6.1550 0.3600 6.3950 0.3600 ;
        POLYGON  3.1950 0.5400 3.0750 0.5400 3.0750 0.5800 2.1350 0.5800 2.1350 1.7300 2.0950 1.7300
                 2.0950 1.8700 1.9750 1.8700 1.9750 1.6100 2.0150 1.6100 2.0150 0.6400 1.8150 0.6400
                 1.8150 0.4000 1.9350 0.4000 1.9350 0.4600 2.9550 0.4600 2.9550 0.4200 3.1950 0.4200 ;
        POLYGON  2.4950 0.8600 2.4850 0.8600 2.4850 2.1100 1.6550 2.1100 1.6550 2.2500 1.4150 2.2500
                 1.4150 2.1300 1.5350 2.1300 1.5350 1.9900 2.3650 1.9900 2.3650 0.8600 2.2550 0.8600
                 2.2550 0.7400 2.4950 0.7400 ;
        POLYGON  1.2950 1.4900 1.0550 1.4900 1.0550 1.7200 0.3950 1.7200 0.3950 1.8100 0.1150 1.8100
                 0.1150 0.5200 0.1350 0.5200 0.1350 0.4000 0.2550 0.4000 0.2550 0.6400 0.2350 0.6400
                 0.2350 1.6000 0.9350 1.6000 0.9350 1.3700 1.2950 1.3700 ;
    END
END DLY3X4

MACRO DLY3X1
    CLASS CORE ;
    FOREIGN DLY3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.4650 2.9250 1.7250 ;
        RECT  2.7050 1.4050 2.9250 1.7250 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3650 1.2300 4.6250 1.3800 ;
        RECT  4.4050 1.1100 4.5250 2.2100 ;
        RECT  4.2650 1.1100 4.5250 1.2300 ;
        RECT  4.2650 0.6800 4.3850 1.2300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  7.1100 1.4800 7.5300 1.7200 ;
        RECT  7.4100 0.9800 7.5300 1.7200 ;
        RECT  7.2050 0.9800 7.5300 1.1000 ;
        RECT  7.2050 -0.1800 7.3250 1.1000 ;
        RECT  6.7250 0.6200 6.8450 0.8600 ;
        RECT  6.6050 -0.1800 6.7250 0.7400 ;
        RECT  5.3250 1.2200 5.5650 1.3400 ;
        RECT  5.4450 -0.1800 5.5650 1.3400 ;
        RECT  4.7450 0.6000 4.9850 0.7200 ;
        RECT  4.8450 -0.1800 4.9650 0.7200 ;
        RECT  3.6350 1.4650 3.8750 1.5850 ;
        RECT  3.6350 -0.1800 3.7550 1.5850 ;
        RECT  2.8350 -0.1800 2.9550 0.8850 ;
        RECT  1.8750 0.7600 1.9950 1.5200 ;
        RECT  1.5750 0.7600 1.9950 0.8800 ;
        RECT  1.5750 -0.1800 1.6950 0.8800 ;
        RECT  1.1750 -0.1800 1.2950 0.6400 ;
        RECT  0.3750 1.3200 0.7950 1.4400 ;
        RECT  0.3750 -0.1800 0.4950 1.4400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  6.1650 1.2200 7.2900 1.3400 ;
        RECT  6.6100 1.9200 6.7300 2.7900 ;
        RECT  6.2300 1.2200 6.3500 2.7900 ;
        RECT  4.7650 1.7000 5.0050 2.1500 ;
        RECT  4.8650 1.7000 4.9850 2.7900 ;
        RECT  3.2750 1.2450 3.5150 1.3650 ;
        RECT  3.2750 1.2450 3.3950 2.7900 ;
        RECT  2.9250 1.8450 3.0450 2.7900 ;
        RECT  0.6150 1.0000 1.7550 1.1200 ;
        RECT  1.1750 1.8900 1.6750 2.0100 ;
        RECT  1.5550 1.0000 1.6750 2.0100 ;
        RECT  1.1750 1.8900 1.4350 2.7900 ;
        RECT  1.0550 1.8000 1.2950 1.9200 ;
        RECT  0.6150 0.7800 0.8550 1.1200 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.7700 1.9800 7.1900 1.9800 7.1900 1.9600 6.8700 1.9600 6.8700 1.6600 6.4700 1.6600
                 6.4700 1.5400 6.9900 1.5400 6.9900 1.8400 7.6500 1.8400 7.6500 0.8600 7.4450 0.8600
                 7.4450 0.6200 7.5650 0.6200 7.5650 0.7400 7.7700 0.7400 ;
        POLYGON  7.0850 1.1000 6.3650 1.1000 6.3650 0.5000 5.8050 0.5000 5.8050 1.5800 5.6450 1.5800
                 5.6450 1.8000 5.5250 1.8000 5.5250 1.4600 5.6850 1.4600 5.6850 0.3800 6.4850 0.3800
                 6.4850 0.9800 6.9650 0.9800 6.9650 0.4800 6.8450 0.4800 6.8450 0.3600 7.0850 0.3600 ;
        POLYGON  6.2450 1.1000 6.0450 1.1000 6.0450 1.9200 6.1100 1.9200 6.1100 2.0400 5.1250 2.0400
                 5.1250 1.5800 4.8650 1.5800 4.8650 1.4200 4.7450 1.4200 4.7450 1.3000 4.9850 1.3000
                 4.9850 1.4600 5.2450 1.4600 5.2450 1.9200 5.9250 1.9200 5.9250 0.9800 6.1250 0.9800
                 6.1250 0.6200 6.2450 0.6200 ;
        POLYGON  5.3250 0.4800 5.2250 0.4800 5.2250 0.9600 4.5050 0.9600 4.5050 0.5600 3.9950 0.5600
                 3.9950 0.7650 4.1150 0.7650 4.1150 1.8250 3.6850 1.8250 3.6850 1.9650 3.5650 1.9650
                 3.5650 1.7050 3.9950 1.7050 3.9950 0.8850 3.8750 0.8850 3.8750 0.4400 4.6250 0.4400
                 4.6250 0.8400 5.1050 0.8400 5.1050 0.4800 5.0850 0.4800 5.0850 0.3600 5.3250 0.3600 ;
        POLYGON  3.3150 0.5050 3.1950 0.5050 3.1950 1.1250 2.5950 1.1250 2.5950 0.5250 2.2350 0.5250
                 2.2350 1.8600 2.1150 1.8600 2.1150 0.6400 1.8150 0.6400 1.8150 0.4000 1.9350 0.4000
                 1.9350 0.4050 2.7150 0.4050 2.7150 1.0050 3.0750 1.0050 3.0750 0.3850 3.3150 0.3850 ;
        POLYGON  2.6250 2.2500 1.5550 2.2500 1.5550 2.1300 2.5050 2.1300 2.5050 1.9650 2.3550 1.9650
                 2.3550 0.6450 2.4750 0.6450 2.4750 1.8450 2.6250 1.8450 ;
        POLYGON  1.4350 1.4800 1.3150 1.4800 1.3150 1.6800 0.5950 1.6800 0.5950 1.8600 0.4750 1.8600
                 0.4750 1.7400 0.1350 1.7400 0.1350 0.4000 0.2550 0.4000 0.2550 1.5600 1.1950 1.5600
                 1.1950 1.3600 1.4350 1.3600 ;
    END
END DLY3X1

MACRO DLY2X4
    CLASS CORE ;
    FOREIGN DLY2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.9600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.6000 1.5150 2.2100 ;
        RECT  1.2150 0.5200 1.5150 0.6400 ;
        RECT  1.3950 0.4000 1.5150 0.6400 ;
        RECT  1.2150 1.6000 1.5150 1.7200 ;
        RECT  1.2150 0.5200 1.3350 1.7200 ;
        RECT  0.5550 0.8850 1.3350 1.0050 ;
        RECT  0.5550 0.8850 0.8000 1.1450 ;
        RECT  0.5550 0.5900 0.6750 2.2100 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 0.7700 3.7000 1.1450 ;
        RECT  3.5050 1.0200 3.6250 1.4000 ;
        END
    END A
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.9600 0.1800 ;
        RECT  6.2400 1.4800 6.6600 1.7200 ;
        RECT  6.5400 0.9800 6.6600 1.7200 ;
        RECT  6.3650 0.9800 6.6600 1.1000 ;
        RECT  6.3650 -0.1800 6.4850 1.1000 ;
        RECT  5.7650 0.6800 6.0050 0.8000 ;
        RECT  5.7650 -0.1800 5.8850 0.8000 ;
        RECT  4.2050 1.3000 4.4850 1.4200 ;
        RECT  4.3650 -0.1800 4.4850 1.4200 ;
        RECT  3.6450 -0.1800 3.8850 0.3200 ;
        RECT  2.4550 1.1000 2.7350 1.2200 ;
        RECT  2.6150 -0.1800 2.7350 1.2200 ;
        RECT  1.8150 -0.1800 1.9350 0.6400 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.9600 2.7900 ;
        RECT  5.2200 1.2200 6.4200 1.3400 ;
        RECT  5.2200 1.8400 5.5800 2.1500 ;
        RECT  5.2200 1.8400 5.4600 2.7900 ;
        RECT  5.2200 1.0600 5.3400 2.7900 ;
        RECT  5.0850 1.0600 5.3400 1.1800 ;
        RECT  3.7250 2.1800 3.8450 2.7900 ;
        RECT  2.2550 0.7600 2.4950 0.9000 ;
        RECT  1.4550 0.7600 2.4950 0.8800 ;
        RECT  1.6350 1.8200 1.9950 2.1500 ;
        RECT  1.6350 1.8200 1.8750 2.7900 ;
        RECT  1.6350 1.3600 1.7550 2.7900 ;
        RECT  1.4550 1.3600 1.7550 1.4800 ;
        RECT  1.4550 0.7600 1.5750 1.4800 ;
        RECT  0.9750 1.5600 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.9000 1.9800 6.3200 1.9800 6.3200 1.9600 6.0000 1.9600 6.0000 1.7200 5.6600 1.7200
                 5.6600 1.4600 5.7800 1.4600 5.7800 1.6000 6.1200 1.6000 6.1200 1.8400 6.7800 1.8400
                 6.7800 0.8600 6.6050 0.8600 6.6050 0.6200 6.7250 0.6200 6.7250 0.7400 6.9000 0.7400 ;
        POLYGON  6.2450 1.0400 5.5250 1.0400 5.5250 0.6200 4.9900 0.6200 4.9900 0.6800 4.7250 0.6800
                 4.7250 1.7000 4.5450 1.7000 4.5450 1.8200 4.4250 1.8200 4.4250 1.5800 4.6050 1.5800
                 4.6050 0.5600 4.8700 0.5600 4.8700 0.5000 5.6450 0.5000 5.6450 0.9200 6.1250 0.9200
                 6.1250 0.4800 6.0050 0.4800 6.0050 0.3600 6.2450 0.3600 ;
        POLYGON  5.4050 0.8600 5.2850 0.8600 5.2850 0.9400 4.9650 0.9400 4.9650 1.5600 5.1000 1.5600
                 5.1000 2.2100 4.9800 2.2100 4.9800 2.0600 3.5600 2.0600 3.5600 2.2200 2.1150 2.2200
                 2.1150 1.7000 1.8750 1.7000 1.8750 1.2400 1.6950 1.2400 1.6950 1.0000 1.8150 1.0000
                 1.8150 1.1200 1.9950 1.1200 1.9950 1.5800 2.2350 1.5800 2.2350 2.1000 3.4400 2.1000
                 3.4400 1.9400 4.8450 1.9400 4.8450 0.8200 5.1650 0.8200 5.1650 0.7400 5.4050 0.7400 ;
        POLYGON  4.2450 0.5400 4.1250 0.5400 4.1250 0.5600 2.9750 0.5600 2.9750 1.4600 2.8350 1.4600
                 2.8350 1.7400 2.5950 1.7400 2.5950 1.6200 2.7150 1.6200 2.7150 1.3400 2.8550 1.3400
                 2.8550 0.4000 2.9750 0.4000 2.9750 0.4400 4.0050 0.4400 4.0050 0.4200 4.2450 0.4200 ;
        POLYGON  3.3650 1.8200 3.3200 1.8200 3.3200 1.9800 2.3550 1.9800 2.3550 1.4600 2.1150 1.4600
                 2.1150 1.2200 2.2350 1.2200 2.2350 1.3400 2.4750 1.3400 2.4750 1.8600 3.2000 1.8600
                 3.2000 1.7000 3.2450 1.7000 3.2450 0.6800 3.3650 0.6800 ;
    END
END DLY2X4

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.8200 2.5400 1.1450 ;
        RECT  2.3300 0.9400 2.4500 1.2600 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2200 1.6000 0.3400 2.1800 ;
        RECT  0.2200 0.4000 0.3400 0.6400 ;
        RECT  0.1000 0.5200 0.2200 1.7200 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.9100 1.4800 5.2100 1.7200 ;
        RECT  5.0900 0.9800 5.2100 1.7200 ;
        RECT  4.9900 -0.1800 5.1100 1.1000 ;
        RECT  4.3900 0.6800 4.6300 0.8000 ;
        RECT  4.3900 -0.1800 4.5100 0.8000 ;
        RECT  3.1900 -0.1800 3.3100 0.7800 ;
        RECT  3.1100 0.6600 3.2300 1.4600 ;
        RECT  2.4700 -0.1800 2.7100 0.3200 ;
        RECT  1.2800 1.0400 1.5600 1.2800 ;
        RECT  1.4400 -0.1800 1.5600 1.2800 ;
        RECT  0.6400 -0.1800 0.7600 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  3.9100 1.2200 4.9700 1.3400 ;
        RECT  4.2900 1.9200 4.5300 2.7900 ;
        RECT  4.2900 1.7000 4.4100 2.7900 ;
        RECT  3.9100 1.7000 4.4100 1.8200 ;
        RECT  3.9100 1.0000 4.0300 1.8200 ;
        RECT  2.4900 2.1800 2.7300 2.3000 ;
        RECT  2.4950 2.1800 2.6150 2.7900 ;
        RECT  1.0800 0.7600 1.3200 0.9000 ;
        RECT  0.3400 0.7600 1.3200 0.8800 ;
        RECT  0.4600 1.8800 0.7600 2.7900 ;
        RECT  0.4600 1.3600 0.5800 2.7900 ;
        RECT  0.3400 0.7600 0.4600 1.4800 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.4500 1.9800 4.9900 1.9800 4.9900 1.9600 4.6700 1.9600 4.6700 1.5800 4.1500 1.5800
                 4.1500 1.4600 4.7900 1.4600 4.7900 1.8400 5.3300 1.8400 5.3300 0.8600 5.2300 0.8600
                 5.2300 0.6200 5.3500 0.6200 5.3500 0.7400 5.4500 0.7400 ;
        POLYGON  4.8700 1.0400 4.1500 1.0400 4.1500 0.5000 3.5500 0.5000 3.5500 1.7000 3.3700 1.7000
                 3.3700 1.8200 3.2500 1.8200 3.2500 1.5800 3.4300 1.5800 3.4300 0.3800 4.2700 0.3800
                 4.2700 0.9200 4.7500 0.9200 4.7500 0.4800 4.6300 0.4800 4.6300 0.3600 4.8700 0.3600 ;
        POLYGON  4.1700 2.0600 2.3700 2.0600 2.3700 2.2500 0.9250 2.2500 0.9250 1.8800 0.8800 1.8800
                 0.8800 1.7600 0.7000 1.7600 0.7000 1.2400 0.5800 1.2400 0.5800 1.0000 0.7000 1.0000
                 0.7000 1.1200 0.8200 1.1200 0.8200 1.6400 1.0000 1.6400 1.0000 1.7600 1.0450 1.7600
                 1.0450 2.1300 2.2500 2.1300 2.2500 1.9400 3.6700 1.9400 3.6700 0.7600 3.9100 0.7600
                 3.9100 0.6200 4.0300 0.6200 4.0300 0.8800 3.7900 0.8800 3.7900 1.9400 4.1700 1.9400 ;
        POLYGON  3.0700 0.5400 2.9500 0.5400 2.9500 0.5600 1.8000 0.5600 1.8000 1.5200 1.5400 1.5200
                 1.5400 1.7700 1.4200 1.7700 1.4200 1.4000 1.6800 1.4000 1.6800 0.4000 1.8000 0.4000
                 1.8000 0.4400 2.8300 0.4400 2.8300 0.4200 3.0700 0.4200 ;
        POLYGON  2.1900 1.8200 2.1300 1.8200 2.1300 2.0100 1.1800 2.0100 1.1800 1.6400 1.1200 1.6400
                 1.1200 1.5200 0.9400 1.5200 0.9400 1.1900 1.0600 1.1900 1.0600 1.4000 1.2400 1.4000
                 1.2400 1.5200 1.3000 1.5200 1.3000 1.8900 2.0100 1.8900 2.0100 1.7000 2.0700 1.7000
                 2.0700 0.6800 2.1900 0.6800 ;
    END
END DLY2X1

MACRO DLY1X4
    CLASS CORE ;
    FOREIGN DLY1X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.0600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.1500 0.5650 1.3800 ;
        RECT  0.3050 1.1500 0.4250 1.5600 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3850 1.3600 3.5050 2.1300 ;
        RECT  2.6800 0.7600 3.5050 0.8800 ;
        RECT  3.3850 0.5900 3.5050 0.8800 ;
        RECT  3.2050 1.3600 3.5050 1.4800 ;
        RECT  2.6800 1.2400 3.3250 1.3600 ;
        RECT  2.6800 1.1750 2.8300 1.4350 ;
        RECT  2.5450 1.3600 2.8000 1.4800 ;
        RECT  2.6800 0.7100 2.8000 1.4800 ;
        RECT  2.5450 0.7100 2.8000 0.8300 ;
        RECT  2.5450 1.3600 2.6650 2.1300 ;
        RECT  2.5450 0.5900 2.6650 0.8300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.0600 0.1800 ;
        RECT  3.8050 -0.1800 3.9250 0.6400 ;
        RECT  2.9650 -0.1800 3.0850 0.6400 ;
        RECT  2.1250 -0.1800 2.2450 0.6400 ;
        RECT  1.1850 1.3600 1.3450 1.6000 ;
        RECT  1.2250 0.7600 1.3450 1.6000 ;
        RECT  0.9550 0.7600 1.3450 0.8800 ;
        RECT  0.9550 -0.1800 1.0750 0.8800 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.0600 2.7900 ;
        RECT  3.8050 1.4800 3.9250 2.7900 ;
        RECT  2.9650 1.4800 3.0850 2.7900 ;
        RECT  2.1250 1.4800 2.2450 2.7900 ;
        RECT  0.9850 1.0000 1.1050 1.2400 ;
        RECT  0.9450 1.1200 1.0650 2.7900 ;
        RECT  0.5550 1.8200 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3850 1.1500 2.2850 1.1500 2.2850 1.3600 1.8250 1.3600 1.8250 2.1300 1.7050 2.1300
                 1.7050 1.2400 2.1650 1.2400 2.1650 0.8800 1.7050 0.8800 1.7050 0.5900 1.8250 0.5900
                 1.8250 0.7600 2.3850 0.7600 ;
        POLYGON  2.0450 1.1200 1.5850 1.1200 1.5850 1.8400 1.3150 1.8400 1.3150 1.9600 1.1950 1.9600
                 1.1950 1.7200 1.4650 1.7200 1.4650 0.6400 1.1950 0.6400 1.1950 0.4000 1.3150 0.4000
                 1.3150 0.5200 1.5850 0.5200 1.5850 1.0000 2.0450 1.0000 ;
        POLYGON  0.8250 1.0300 0.1850 1.0300 0.1850 1.6800 0.2550 1.6800 0.2550 1.9400 0.1350 1.9400
                 0.1350 1.8000 0.0650 1.8000 0.0650 0.5200 0.1350 0.5200 0.1350 0.4000 0.2550 0.4000
                 0.2550 0.6400 0.1850 0.6400 0.1850 0.9100 0.8250 0.9100 ;
    END
END DLY1X4

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5300 1.1750 0.8000 1.4350 ;
        RECT  0.3950 1.1800 0.8000 1.4200 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7350 0.6700 2.8550 2.2100 ;
        RECT  2.6800 0.8850 2.8550 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.3150 -0.1800 2.4350 0.7200 ;
        RECT  1.1950 1.3200 1.4750 1.4400 ;
        RECT  1.3550 0.7600 1.4750 1.4400 ;
        RECT  0.9550 0.7600 1.4750 0.8800 ;
        RECT  0.9550 -0.1800 1.0750 0.8800 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.3150 1.5600 2.4350 2.7900 ;
        RECT  0.9550 1.0000 1.2350 1.1200 ;
        RECT  0.9550 1.0000 1.0750 2.7900 ;
        RECT  0.5550 1.7000 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.5600 1.2300 2.4150 1.2300 2.4150 1.4400 1.9550 1.4400 1.9550 1.8000 1.8350 1.8000
                 1.8350 1.3200 2.2950 1.3200 2.2950 0.9600 1.8350 0.9600 1.8350 0.6700 1.9550 0.6700
                 1.9550 0.8400 2.5600 0.8400 ;
        POLYGON  2.1750 1.2000 1.7150 1.2000 1.7150 1.6800 1.3150 1.6800 1.3150 1.8200 1.1950 1.8200
                 1.1950 1.5600 1.5950 1.5600 1.5950 0.6400 1.1950 0.6400 1.1950 0.4000 1.3150 0.4000
                 1.3150 0.5200 1.7150 0.5200 1.7150 1.0800 2.1750 1.0800 ;
        POLYGON  0.8350 1.0000 0.2550 1.0000 0.2550 1.8200 0.1350 1.8200 0.1350 0.4000 0.2550 0.4000
                 0.2550 0.8800 0.8350 0.8800 ;
    END
END DLY1X1

MACRO DFFXL
    CLASS CORE ;
    FOREIGN DFFXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0300 1.1550 2.3050 1.3800 ;
        RECT  1.9250 1.1200 2.1850 1.3150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3950 1.4800 6.6950 1.7300 ;
        RECT  6.3950 1.4800 6.6550 1.7500 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 1.3000 0.2550 1.5800 ;
        RECT  0.1350 0.6800 0.2550 0.9400 ;
        RECT  0.1150 0.8200 0.2350 1.4200 ;
        RECT  0.0700 0.8850 0.2350 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.3800 1.5650 1.6200 ;
        RECT  1.3650 0.6800 1.4850 0.9600 ;
        RECT  1.3250 0.8400 1.4450 1.6200 ;
        RECT  1.2300 1.4650 1.3800 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.5150 0.6700 6.7550 0.7900 ;
        RECT  6.6350 -0.1800 6.7550 0.7900 ;
        RECT  5.0150 0.5700 5.2550 0.6900 ;
        RECT  5.1350 -0.1800 5.2550 0.6900 ;
        RECT  3.0950 -0.1800 3.2150 0.8600 ;
        RECT  1.8050 -0.1800 1.9250 0.4000 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.5950 1.8700 6.7150 2.7900 ;
        RECT  4.9550 2.2900 5.1950 2.7900 ;
        RECT  3.1750 2.2900 3.4150 2.7900 ;
        RECT  1.8650 1.5000 1.9850 2.7900 ;
        RECT  0.5550 1.4600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.1750 1.5100 7.1350 1.5100 7.1350 1.9900 7.0150 1.9900 7.0150 1.3900 7.0550 1.3900
                 7.0550 1.0300 6.2750 1.0300 6.2750 0.5000 5.5950 0.5000 5.5950 0.9300 4.7750 0.9300
                 4.7750 0.5000 4.4150 0.5000 4.4150 1.1200 4.2950 1.1200 4.2950 1.3300 3.7750 1.3300
                 3.7750 1.4500 3.6550 1.4500 3.6550 1.2100 4.1750 1.2100 4.1750 1.0000 4.2950 1.0000
                 4.2950 0.3800 4.8950 0.3800 4.8950 0.8100 5.4750 0.8100 5.4750 0.3800 5.5750 0.3800
                 5.5750 0.3600 5.8150 0.3600 5.8150 0.3800 6.3950 0.3800 6.3950 0.9100 7.0550 0.9100
                 7.0550 0.6200 7.1750 0.6200 ;
        POLYGON  6.9350 1.2700 6.8150 1.2700 6.8150 1.3600 6.2750 1.3600 6.2750 1.4000 6.0750 1.4000
                 6.0750 2.2300 5.3150 2.2300 5.3150 2.1700 4.3550 2.1700 4.3550 2.2300 3.6100 2.2300
                 3.6100 2.1700 2.2850 2.1700 2.2850 1.5000 2.4250 1.5000 2.4250 1.0000 2.2850 1.0000
                 2.2850 0.6800 2.4050 0.6800 2.4050 0.8800 2.5450 0.8800 2.5450 1.6200 2.4050 1.6200
                 2.4050 2.0500 3.7300 2.0500 3.7300 2.1100 4.2350 2.1100 4.2350 1.6100 4.1750 1.6100
                 4.1750 1.4900 4.4150 1.4900 4.4150 1.6100 4.3550 1.6100 4.3550 2.0500 5.4350 2.0500
                 5.4350 2.1100 5.9550 2.1100 5.9550 1.6100 5.5150 1.6100 5.5150 1.4900 5.9550 1.4900
                 5.9550 1.2400 6.1550 1.2400 6.1550 1.1600 6.2750 1.1600 6.2750 1.2400 6.6950 1.2400
                 6.6950 1.1500 6.9350 1.1500 ;
        POLYGON  5.9950 0.8600 5.8350 0.8600 5.8350 1.3700 5.3950 1.3700 5.3950 1.7300 5.8350 1.7300
                 5.8350 1.9900 5.7150 1.9900 5.7150 1.8500 5.2750 1.8500 5.2750 1.5300 4.9150 1.5300
                 4.9150 1.6500 4.7950 1.6500 4.7950 1.4100 5.2750 1.4100 5.2750 1.2500 5.7150 1.2500
                 5.7150 0.7400 5.8750 0.7400 5.8750 0.6200 5.9950 0.6200 ;
        POLYGON  5.1550 1.2900 4.6550 1.2900 4.6550 1.8100 4.7150 1.8100 4.7150 1.9300 4.4750 1.9300
                 4.4750 1.8100 4.5350 1.8100 4.5350 0.6200 4.6550 0.6200 4.6550 1.1700 5.0350 1.1700
                 5.0350 1.0500 5.1550 1.0500 ;
        POLYGON  4.1750 0.8000 3.7900 0.8000 3.7900 1.0900 3.5350 1.0900 3.5350 1.5700 4.0550 1.5700
                 4.0550 1.9900 3.9350 1.9900 3.9350 1.6900 3.4150 1.6900 3.4150 1.6500 3.0150 1.6500
                 3.0150 1.4100 3.1350 1.4100 3.1350 1.5300 3.4150 1.5300 3.4150 0.9700 3.6700 0.9700
                 3.6700 0.6800 4.1750 0.6800 ;
        POLYGON  3.2950 1.2200 2.8950 1.2200 2.8950 1.8100 2.9350 1.8100 2.9350 1.9300 2.6950 1.9300
                 2.6950 1.8100 2.7750 1.8100 2.7750 0.8600 2.6750 0.8600 2.6750 0.5600 2.1650 0.5600
                 2.1650 1.0000 1.8050 1.0000 1.8050 1.2000 1.5650 1.2000 1.5650 1.0800 1.6850 1.0800
                 1.6850 0.8800 2.0450 0.8800 2.0450 0.4400 2.7950 0.4400 2.7950 0.7400 2.8950 0.7400
                 2.8950 1.1000 3.1750 1.1000 3.1750 0.9800 3.2950 0.9800 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.1800 0.3550 1.1800 0.3550 1.0600 0.9750 1.0600
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFXL

MACRO DFFX4
    CLASS CORE ;
    FOREIGN DFFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.8850 0.3950 1.1250 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5450 1.3150 1.6650 1.5550 ;
        RECT  1.2300 1.3150 1.6650 1.4350 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7050 0.7200 6.9050 0.8400 ;
        RECT  6.7650 1.4400 6.8850 2.2100 ;
        RECT  6.5850 1.4400 6.8850 1.5600 ;
        RECT  5.9000 1.3200 6.7050 1.4400 ;
        RECT  5.9250 0.7200 6.0450 2.2100 ;
        RECT  5.8700 1.1750 6.0450 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6250 0.7200 8.8250 0.8400 ;
        RECT  8.4450 1.4400 8.5650 2.2100 ;
        RECT  8.2650 1.4400 8.5650 1.5600 ;
        RECT  7.6100 1.3200 8.3850 1.4400 ;
        RECT  7.6400 0.7200 7.7600 1.5600 ;
        RECT  7.6050 1.4400 7.7250 2.2100 ;
        RECT  7.6100 1.1750 7.7600 1.5600 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.1850 -0.1800 9.3050 0.7100 ;
        RECT  8.1050 -0.1800 8.3450 0.3600 ;
        RECT  7.1450 -0.1800 7.3850 0.3600 ;
        RECT  6.1850 -0.1800 6.4250 0.3600 ;
        RECT  5.2250 -0.1800 5.4650 0.3600 ;
        RECT  4.3250 -0.1800 4.4450 0.3800 ;
        RECT  2.7250 -0.1800 2.8450 0.3800 ;
        RECT  1.4850 -0.1800 1.6050 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  8.8650 1.5800 8.9850 2.7900 ;
        RECT  8.0250 1.5600 8.1450 2.7900 ;
        RECT  7.1850 1.5600 7.3050 2.7900 ;
        RECT  6.3450 1.5600 6.4650 2.7900 ;
        RECT  5.5050 1.5600 5.6250 2.7900 ;
        RECT  4.6050 1.6700 4.7250 2.7900 ;
        RECT  2.8250 2.2600 3.0650 2.7900 ;
        RECT  1.3850 1.9500 1.5050 2.7900 ;
        RECT  0.1350 1.4600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.7250 0.9000 9.5450 0.9000 9.5450 1.4600 9.4050 1.4600 9.4050 2.2100 9.2850 2.2100
                 9.2850 1.4600 8.7250 1.4600 8.7250 1.2200 8.8450 1.2200 8.8450 1.3400 9.4250 1.3400
                 9.4250 0.7800 9.6050 0.7800 9.6050 0.6600 9.7250 0.6600 ;
        POLYGON  9.2650 1.2200 9.1450 1.2200 9.1450 0.9500 8.9450 0.9500 8.9450 0.6000 5.1650 0.6000
                 5.1650 1.3200 5.6300 1.3200 5.6300 1.2000 5.7500 1.2000 5.7500 1.4400 5.1450 1.4400
                 5.1450 2.1900 5.0250 2.1900 5.0250 1.4400 4.6850 1.4400 4.6850 1.5000 4.4450 1.5000
                 4.4450 1.3800 4.5650 1.3800 4.5650 1.3200 5.0450 1.3200 5.0450 0.8000 4.8050 0.8000
                 4.8050 0.5600 4.9250 0.5600 4.9250 0.6800 5.0450 0.6800 5.0450 0.4800 9.0650 0.4800
                 9.0650 0.8300 9.2650 0.8300 ;
        POLYGON  4.9250 1.1600 3.9450 1.1600 3.9450 1.8900 4.0850 1.8900 4.0850 2.0100 3.8250 2.0100
                 3.8250 0.8400 3.6850 0.8400 3.6850 0.7200 3.9450 0.7200 3.9450 1.0400 4.9250 1.0400 ;
        POLYGON  4.3250 2.2500 3.1850 2.2500 3.1850 2.1400 2.7050 2.1400 2.7050 2.2500 1.8650 2.2500
                 1.8650 1.7950 1.1100 1.7950 1.1100 1.9150 1.0850 1.9150 1.0850 2.0700 0.9650 2.0700
                 0.9650 1.7950 0.9900 1.7950 0.9900 0.8400 0.8850 0.8400 0.8850 0.7200 1.1250 0.7200
                 1.1250 0.8400 1.1100 0.8400 1.1100 1.6750 1.8650 1.6750 1.8650 1.4900 1.9850 1.4900
                 1.9850 2.1300 2.5850 2.1300 2.5850 2.0200 3.3050 2.0200 3.3050 2.1300 4.2050 2.1300
                 4.2050 1.7300 4.0650 1.7300 4.0650 1.4900 4.1850 1.4900 4.1850 1.6100 4.3250 1.6100 ;
        POLYGON  4.0850 0.5000 3.9650 0.5000 3.9650 0.5400 3.5650 0.5400 3.5650 1.4200 3.7050 1.4200
                 3.7050 1.6600 3.5850 1.6600 3.5850 1.5400 3.4450 1.5400 3.4450 0.5400 3.0850 0.5400
                 3.0850 0.6200 2.4650 0.6200 2.4650 1.6600 2.3450 1.6600 2.3450 0.6000 1.8450 0.6000
                 1.8450 0.6200 1.2450 0.6200 1.2450 0.6000 0.6750 0.6000 0.6750 1.5800 0.5550 1.5800
                 0.5550 0.4800 1.0450 0.4800 1.0450 0.3800 1.3650 0.3800 1.3650 0.5000 1.7250 0.5000
                 1.7250 0.4800 1.8050 0.4800 1.8050 0.3800 2.0450 0.3800 2.0450 0.4800 2.4650 0.4800
                 2.4650 0.5000 2.9650 0.5000 2.9650 0.4200 3.8450 0.4200 3.8450 0.3800 4.0850 0.3800 ;
        POLYGON  3.6650 2.0100 3.4250 2.0100 3.4250 1.9000 3.2050 1.9000 3.2050 1.3200 2.6850 1.3200
                 2.6850 1.0800 2.8050 1.0800 2.8050 1.2000 3.2050 1.2000 3.2050 0.6600 3.3250 0.6600
                 3.3250 1.7800 3.5450 1.7800 3.5450 1.8900 3.6650 1.8900 ;
        POLYGON  3.0850 1.6900 2.9650 1.6900 2.9650 1.9000 2.3450 1.9000 2.3450 2.0100 2.1050 2.0100
                 2.1050 0.8400 1.9650 0.8400 1.9650 0.7200 2.2250 0.7200 2.2250 1.7800 2.8450 1.7800
                 2.8450 1.5700 3.0850 1.5700 ;
    END
END DFFX4

MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8150 1.3100 0.9350 1.5500 ;
        RECT  0.5950 1.5200 0.8550 1.6700 ;
        RECT  0.7350 1.4300 0.9350 1.5500 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 0.8050 5.1500 1.1450 ;
        RECT  4.9550 0.9200 5.0750 1.2600 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5800 0.8850 5.7300 1.1450 ;
        RECT  5.5950 0.6800 5.7150 2.0300 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5550 0.6800 6.6750 0.9700 ;
        RECT  6.4350 0.8500 6.5550 2.0300 ;
        RECT  6.1600 0.9700 6.5550 1.0900 ;
        RECT  6.1600 0.8850 6.3100 1.1450 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  7.0350 -0.1800 7.1550 0.7300 ;
        RECT  6.0150 -0.1800 6.2550 0.3200 ;
        RECT  5.0550 -0.1800 5.2950 0.3200 ;
        RECT  3.7350 -0.1800 3.8550 0.8200 ;
        RECT  2.1150 -0.1800 2.3550 0.3200 ;
        RECT  0.6750 -0.1800 0.7950 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  6.8550 1.3800 6.9750 2.7900 ;
        RECT  6.0150 1.3800 6.1350 2.7900 ;
        RECT  5.1750 1.3800 5.2950 2.7900 ;
        RECT  3.7550 2.1300 3.9950 2.2500 ;
        RECT  3.7550 2.1300 3.8750 2.7900 ;
        RECT  2.0150 2.1700 2.2550 2.2900 ;
        RECT  2.0150 2.1700 2.1350 2.7900 ;
        RECT  0.6150 1.7900 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.7550 0.8600 7.6350 0.8600 7.6350 1.2100 7.4550 1.2100 7.4550 1.6200 7.3350 1.6200
                 7.3350 1.2100 6.6750 1.2100 6.6750 1.0900 7.5150 1.0900 7.5150 0.7400 7.7550 0.7400 ;
        POLYGON  7.5350 0.5200 7.3950 0.5200 7.3950 0.9700 6.7950 0.9700 6.7950 0.5600 5.9950 0.5600
                 5.9950 1.2400 5.8750 1.2400 5.8750 0.5600 5.4350 0.5600 5.4350 1.2400 5.3150 1.2400
                 5.3150 0.5600 4.2750 0.5600 4.2750 0.8000 4.5550 0.8000 4.5550 1.4500 4.4750 1.4500
                 4.4750 1.7700 4.2350 1.7700 4.2350 1.6500 4.3550 1.6500 4.3550 1.4500 3.7350 1.4500
                 3.7350 1.3300 4.4350 1.3300 4.4350 0.9200 4.1550 0.9200 4.1550 0.4400 6.9150 0.4400
                 6.9150 0.8500 7.2750 0.8500 7.2750 0.4000 7.5350 0.4000 ;
        POLYGON  4.8150 2.0100 3.5350 2.0100 3.5350 2.0500 3.0750 2.0500 3.0750 2.2500 2.8350 2.2500
                 2.8350 2.0500 1.8950 2.0500 1.8950 2.2500 1.4550 2.2500 1.4550 2.1300 1.7750 2.1300
                 1.7750 1.9300 3.4150 1.9300 3.4150 1.8900 4.6950 1.8900 4.6950 1.6200 4.6750 1.6200
                 4.6750 0.6800 4.7950 0.6800 4.7950 1.5000 4.8150 1.5000 ;
        POLYGON  4.3150 1.2000 4.0750 1.2000 4.0750 1.1700 3.6150 1.1700 3.6150 1.7700 3.2950 1.7700
                 3.2950 1.8100 3.0550 1.8100 3.0550 1.6900 3.1750 1.6900 3.1750 1.6500 3.4950 1.6500
                 3.4950 1.1700 3.0350 1.1700 3.0350 0.6800 3.1550 0.6800 3.1550 1.0500 4.1950 1.0500
                 4.1950 1.0800 4.3150 1.0800 ;
        POLYGON  3.3750 1.5300 3.2550 1.5300 3.2550 1.4100 2.7950 1.4100 2.7950 1.2800 2.7150 1.2800
                 2.7150 1.0400 2.7950 1.0400 2.7950 0.5600 1.2350 0.5600 1.2350 1.3700 1.3550 1.3700
                 1.3550 1.4900 1.1150 1.4900 1.1150 1.1600 0.3750 1.1600 0.3750 1.7500 0.2550 1.7500
                 0.2550 1.8700 0.1350 1.8700 0.1350 1.6300 0.2550 1.6300 0.2550 0.6800 0.3750 0.6800
                 0.3750 1.0400 1.1150 1.0400 1.1150 0.4400 1.5550 0.4400 1.5550 0.4200 1.7950 0.4200
                 1.7950 0.4400 2.9150 0.4400 2.9150 1.2900 3.3750 1.2900 ;
        POLYGON  2.7350 1.8100 2.4950 1.8100 2.4950 1.5200 1.8950 1.5200 1.8950 1.4900 1.7750 1.4900
                 1.7750 1.3700 2.0150 1.3700 2.0150 1.4000 2.4750 1.4000 2.4750 0.8000 2.5550 0.8000
                 2.5550 0.6800 2.6750 0.6800 2.6750 0.9200 2.5950 0.9200 2.5950 1.4000 2.6150 1.4000
                 2.6150 1.6900 2.7350 1.6900 ;
        POLYGON  2.3550 1.2500 1.5950 1.2500 1.5950 1.7500 1.4350 1.7500 1.4350 1.8700 1.3150 1.8700
                 1.3150 1.6300 1.4750 1.6300 1.4750 0.6800 1.5950 0.6800 1.5950 1.1300 2.3550 1.1300 ;
    END
END DFFX2

MACRO DFFX1
    CLASS CORE ;
    FOREIGN DFFX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.2500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8600 1.2100 2.1400 1.3300 ;
        RECT  2.0200 1.0900 2.1400 1.3300 ;
        RECT  1.8100 1.4650 1.9800 1.7250 ;
        RECT  1.8600 1.2100 1.9800 1.7250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3950 1.4500 6.6550 1.6700 ;
        RECT  6.4350 1.3600 6.5550 1.7500 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3800 0.6800 1.5000 2.0800 ;
        RECT  1.2300 0.8850 1.5000 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.2500 0.1800 ;
        RECT  6.5150 -0.1800 6.6350 0.7600 ;
        RECT  4.9550 0.3500 5.1950 0.4700 ;
        RECT  4.9550 -0.1800 5.0750 0.4700 ;
        RECT  3.2350 -0.1800 3.3550 0.8600 ;
        RECT  1.8000 -0.1800 1.9200 0.7300 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.2500 2.7900 ;
        RECT  6.4950 1.8700 6.6150 2.7900 ;
        RECT  4.8950 2.2900 5.1350 2.7900 ;
        RECT  3.1150 2.2900 3.3550 2.7900 ;
        RECT  1.8600 2.0700 1.9800 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.1750 1.4800 7.0350 1.4800 7.0350 1.9900 6.9150 1.9900 6.9150 1.3600 7.0550 1.3600
                 7.0550 0.8600 6.9250 0.8600 6.9250 1.0000 6.2750 1.0000 6.2750 0.5000 5.4350 0.5000
                 5.4350 0.7100 4.7150 0.7100 4.7150 0.5000 4.3550 0.5000 4.3550 1.0700 4.4350 1.0700
                 4.4350 1.3100 4.3150 1.3100 4.3150 1.1900 3.8950 1.1900 3.8950 1.6500 3.7750 1.6500
                 3.7750 1.0700 4.2350 1.0700 4.2350 0.3800 4.8350 0.3800 4.8350 0.5900 5.3150 0.5900
                 5.3150 0.3800 5.5150 0.3800 5.5150 0.3600 5.7550 0.3600 5.7550 0.3800 6.3950 0.3800
                 6.3950 0.8800 6.8050 0.8800 6.8050 0.7400 6.9950 0.7400 6.9950 0.6200 7.1150 0.6200
                 7.1150 0.7400 7.1750 0.7400 ;
        POLYGON  6.9350 1.2400 6.2750 1.2400 6.2750 1.3400 6.0750 1.3400 6.0750 2.1700 2.3050 2.1700
                 2.3050 1.5500 2.2800 1.5500 2.2800 0.6800 2.4000 0.6800 2.4000 1.4300 2.4250 1.4300
                 2.4250 2.0500 4.1750 2.0500 4.1750 1.6700 4.1550 1.6700 4.1550 1.4300 4.2750 1.4300
                 4.2750 1.5500 4.2950 1.5500 4.2950 2.0500 5.9550 2.0500 5.9550 1.6700 5.5150 1.6700
                 5.5150 1.4300 5.6350 1.4300 5.6350 1.5500 5.9550 1.5500 5.9550 1.1200 6.9350 1.1200 ;
        POLYGON  5.9350 1.0000 5.8350 1.0000 5.8350 1.3100 5.3950 1.3100 5.3950 1.7900 5.7150 1.7900
                 5.7150 1.8100 5.8350 1.8100 5.8350 1.9300 5.5950 1.9300 5.5950 1.9100 5.2750 1.9100
                 5.2750 1.5500 4.9150 1.5500 4.9150 1.6700 4.7950 1.6700 4.7950 1.4300 5.2750 1.4300
                 5.2750 1.1900 5.7150 1.1900 5.7150 0.8800 5.8150 0.8800 5.8150 0.6200 5.9350 0.6200 ;
        POLYGON  5.1550 1.2900 4.6750 1.2900 4.6750 1.9300 4.4150 1.9300 4.4150 1.8100 4.5550 1.8100
                 4.5550 0.9500 4.4750 0.9500 4.4750 0.6200 4.5950 0.6200 4.5950 0.8300 4.6750 0.8300
                 4.6750 1.1700 5.1550 1.1700 ;
        POLYGON  4.1150 0.8000 3.6550 0.8000 3.6550 1.7700 3.9350 1.7700 3.9350 1.8100 4.0550 1.8100
                 4.0550 1.9300 3.8150 1.9300 3.8150 1.8900 3.5350 1.8900 3.5350 1.6700 2.9350 1.6700
                 2.9350 1.4300 3.0550 1.4300 3.0550 1.5500 3.5350 1.5500 3.5350 0.6800 4.1150 0.6800 ;
        POLYGON  3.4150 1.4300 3.2950 1.4300 3.2950 1.3100 2.8150 1.3100 2.8150 1.8100 2.8750 1.8100
                 2.8750 1.9300 2.6350 1.9300 2.6350 1.8100 2.6950 1.8100 2.6950 0.7400 2.7950 0.7400
                 2.7950 0.5600 2.1600 0.5600 2.1600 0.9700 1.7400 0.9700 1.7400 1.2400 1.6200 1.2400
                 1.6200 0.8500 2.0400 0.8500 2.0400 0.4400 2.9150 0.4400 2.9150 0.8600 2.8150 0.8600
                 2.8150 1.1900 3.4150 1.1900 ;
        POLYGON  1.1100 1.5800 0.9900 1.5800 0.9900 1.2000 0.3750 1.2000 0.3750 1.0800 0.9900 1.0800
                 0.9900 0.6800 1.1100 0.6800 ;
    END
END DFFX1

MACRO DFFTRXL
    CLASS CORE ;
    FOREIGN DFFTRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9650 1.2700 2.0850 1.5100 ;
        RECT  1.8400 1.3900 2.0850 1.5100 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7400 1.0250 7.0950 1.1600 ;
        RECT  6.7400 0.8850 6.8900 1.1800 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3350 0.7350 7.4550 1.2400 ;
        RECT  7.0300 0.7350 7.4550 0.8550 ;
        RECT  7.0300 0.5950 7.1800 0.8550 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 1.3100 1.4850 1.8300 ;
        RECT  1.3650 0.6700 1.4850 0.9100 ;
        RECT  1.2300 1.1750 1.4450 1.4350 ;
        RECT  1.3250 0.7900 1.4450 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  6.8650 -0.1800 6.9850 0.3800 ;
        RECT  4.7300 -0.1800 4.9700 0.3200 ;
        RECT  3.1350 -0.1800 3.2550 0.9000 ;
        RECT  1.7850 -0.1800 1.9050 0.3900 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  7.5750 1.9800 7.6950 2.7900 ;
        RECT  6.8350 1.9800 6.9550 2.7900 ;
        RECT  4.7150 2.1600 4.9550 2.2800 ;
        RECT  4.7150 2.1600 4.8350 2.7900 ;
        RECT  3.0150 2.1600 3.2550 2.2800 ;
        RECT  3.0150 2.1600 3.1350 2.7900 ;
        RECT  1.7250 2.2300 1.8450 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.6950 1.4800 7.3150 1.4800 7.3150 1.7600 6.0150 1.7600 6.0150 1.8600 5.8950 1.8600
                 5.8950 1.6200 6.0550 1.6200 6.0550 0.9000 5.9950 0.9000 5.9950 0.6600 6.1150 0.6600
                 6.1150 0.7800 6.1750 0.7800 6.1750 1.6400 7.1950 1.6400 7.1950 1.3600 7.5750 1.3600
                 7.5750 0.6600 7.6950 0.6600 ;
        POLYGON  6.5350 1.5200 6.2950 1.5200 6.2950 1.4000 6.3850 1.4000 6.3850 0.6600 6.2850 0.6600
                 6.2850 0.5400 5.8750 0.5400 5.8750 1.3600 5.9350 1.3600 5.9350 1.4800 5.6950 1.4800
                 5.6950 1.3600 5.7550 1.3600 5.7550 0.5400 5.2100 0.5400 5.2100 0.5600 4.1750 0.5600
                 4.1750 1.0000 4.3150 1.0000 4.3150 1.2400 4.0550 1.2400 4.0550 1.1400 3.7550 1.1400
                 3.7550 1.5400 3.6350 1.5400 3.6350 1.0200 4.0550 1.0200 4.0550 0.4400 5.0900 0.4400
                 5.0900 0.4200 5.2350 0.4200 5.2350 0.3800 5.4750 0.3800 5.4750 0.4200 6.4050 0.4200
                 6.4050 0.5400 6.5050 0.5400 6.5050 1.4000 6.5350 1.4000 ;
        POLYGON  5.6350 0.8400 5.5750 0.8400 5.5750 1.6200 5.5950 1.6200 5.5950 1.8600 5.4750 1.8600
                 5.4750 1.7400 5.4550 1.7400 5.4550 1.4800 4.6750 1.4800 4.6750 1.3600 5.4550 1.3600
                 5.4550 0.8400 5.3950 0.8400 5.3950 0.7200 5.6350 0.7200 ;
        POLYGON  5.5150 2.2400 5.2750 2.2400 5.2750 2.1000 5.1750 2.1000 5.1750 2.0400 4.2350 2.0400
                 4.2350 2.2400 3.9950 2.2400 3.9950 2.0400 2.2050 2.0400 2.2050 1.6800 2.2650 1.6800
                 2.2650 0.6700 2.3850 0.6700 2.3850 1.8000 2.3250 1.8000 2.3250 1.9200 5.2950 1.9200
                 5.2950 1.9800 5.3950 1.9800 5.3950 2.1200 5.5150 2.1200 ;
        POLYGON  5.1350 1.1600 4.5550 1.1600 4.5550 1.8000 4.2350 1.8000 4.2350 1.6800 4.4350 1.6800
                 4.4350 0.8400 4.2950 0.8400 4.2950 0.7200 4.5550 0.7200 4.5550 1.0400 5.1350 1.0400 ;
        POLYGON  3.9550 1.8000 3.7150 1.8000 3.7150 1.7800 3.3950 1.7800 3.3950 1.5000 2.9150 1.5000
                 2.9150 1.4600 2.7550 1.4600 2.7550 1.3400 3.0350 1.3400 3.0350 1.3800 3.3950 1.3800
                 3.3950 0.7800 3.8150 0.7800 3.8150 0.6600 3.9350 0.6600 3.9350 0.9000 3.5150 0.9000
                 3.5150 1.6600 3.8350 1.6600 3.8350 1.6800 3.9550 1.6800 ;
        POLYGON  3.2750 1.2600 3.1550 1.2600 3.1550 1.2200 2.6350 1.2200 2.6350 1.6800 2.7750 1.6800
                 2.7750 1.8000 2.5150 1.8000 2.5150 0.7800 2.6550 0.7800 2.6550 0.6600 2.5550 0.6600
                 2.5550 0.5500 2.1450 0.5500 2.1450 1.1500 1.8050 1.1500 1.8050 1.1900 1.5650 1.1900
                 1.5650 1.0300 2.0250 1.0300 2.0250 0.4300 2.6750 0.4300 2.6750 0.5400 2.7750 0.5400
                 2.7750 0.9000 2.6350 0.9000 2.6350 1.1000 3.1550 1.1000 3.1550 1.0200 3.2750 1.0200 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFTRXL

MACRO DFFTRX4
    CLASS CORE ;
    FOREIGN DFFTRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.7300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1650 1.1000 0.3550 1.3400 ;
        RECT  0.0700 1.1750 0.2850 1.4350 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6400 1.1000 0.8000 1.5250 ;
        RECT  0.6650 1.0800 0.7950 1.5250 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.1850 1.7250 1.3800 ;
        RECT  1.4650 1.0200 1.5850 1.3800 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5750 0.7400 7.7750 0.8600 ;
        RECT  7.6350 1.4400 7.7550 2.2100 ;
        RECT  7.4550 1.4400 7.7550 1.5600 ;
        RECT  6.7700 1.3200 7.5750 1.4400 ;
        RECT  6.7950 0.7400 6.9150 2.2100 ;
        RECT  6.7400 1.1750 6.9150 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4950 0.7400 9.6950 0.8600 ;
        RECT  9.3150 1.3200 9.4350 2.2100 ;
        RECT  8.4800 1.3200 9.4350 1.4400 ;
        RECT  8.5100 0.7400 8.6300 1.5600 ;
        RECT  8.4750 1.4400 8.5950 2.2100 ;
        RECT  8.4800 1.1750 8.6300 1.5600 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.7300 0.1800 ;
        RECT  10.0550 -0.1800 10.1750 0.7300 ;
        RECT  8.9750 -0.1800 9.2150 0.3800 ;
        RECT  8.0150 -0.1800 8.2550 0.3800 ;
        RECT  7.0550 -0.1800 7.2950 0.3800 ;
        RECT  6.0950 -0.1800 6.3350 0.3800 ;
        RECT  5.2550 -0.1800 5.3750 0.9200 ;
        RECT  3.6050 -0.1800 3.8450 0.3200 ;
        RECT  1.6150 -0.1800 1.7350 0.6600 ;
        RECT  0.1650 -0.1800 0.2850 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.7300 2.7900 ;
        RECT  9.7350 1.6000 9.8550 2.7900 ;
        RECT  8.8950 1.5600 9.0150 2.7900 ;
        RECT  8.0550 1.5600 8.1750 2.7900 ;
        RECT  7.2150 1.5600 7.3350 2.7900 ;
        RECT  6.3750 1.5600 6.4950 2.7900 ;
        RECT  5.4750 1.6400 5.5950 2.7900 ;
        RECT  3.6050 1.7500 3.7250 2.7900 ;
        RECT  1.7650 1.9800 1.8850 2.7900 ;
        RECT  0.9750 1.9800 1.0950 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.5950 0.9200 10.4150 0.9200 10.4150 1.4800 10.2750 1.4800 10.2750 2.2100
                 10.1550 2.2100 10.1550 1.4800 9.5550 1.4800 9.5550 1.3000 9.7950 1.3000 9.7950 1.3600
                 10.2950 1.3600 10.2950 0.8000 10.4750 0.8000 10.4750 0.6800 10.5950 0.6800 ;
        POLYGON  10.1350 1.2400 10.0150 1.2400 10.0150 0.9700 9.8150 0.9700 9.8150 0.6200 6.3250 0.6200
                 6.3250 0.6800 5.7950 0.6800 5.7950 0.8000 6.1550 0.8000 6.1550 1.3000 6.6200 1.3000
                 6.6200 1.4200 6.0150 1.4200 6.0150 2.1500 5.8950 2.1500 5.8950 1.4200 5.5150 1.4200
                 5.5150 1.5200 5.3950 1.5200 5.3950 1.2800 5.5150 1.2800 5.5150 1.3000 6.0350 1.3000
                 6.0350 0.9200 5.6750 0.9200 5.6750 0.5600 6.2050 0.5600 6.2050 0.5000 9.9350 0.5000
                 9.9350 0.8500 10.1350 0.8500 ;
        POLYGON  5.9150 1.1800 5.6750 1.1800 5.6750 1.1600 5.2750 1.1600 5.2750 1.7700 4.9350 1.7700
                 4.9350 1.8100 4.6950 1.8100 4.6950 1.6900 4.8150 1.6900 4.8150 1.6500 5.1550 1.6500
                 5.1550 1.1600 4.6150 1.1600 4.6150 0.6800 4.7350 0.6800 4.7350 1.0400 5.9150 1.0400 ;
        POLYGON  5.0350 1.5300 4.9150 1.5300 4.9150 1.4000 4.3750 1.4000 4.3750 0.5600 2.7850 0.5600
                 2.7850 1.3700 2.8450 1.3700 2.8450 1.4900 2.6050 1.4900 2.6050 1.3700 2.6650 1.3700
                 2.6650 0.5600 2.2450 0.5600 2.2450 1.5800 2.1250 1.5800 2.1250 0.6600 2.0350 0.6600
                 2.0350 0.4200 2.1550 0.4200 2.1550 0.4400 3.0650 0.4400 3.0650 0.4000 3.3050 0.4000
                 3.3050 0.4400 4.4950 0.4400 4.4950 1.2800 5.0350 1.2800 ;
        POLYGON  4.2550 1.8700 4.1350 1.8700 4.1350 1.4900 3.4050 1.4900 3.4050 1.3700 4.1350 1.3700
                 4.1350 0.6800 4.2550 0.6800 ;
        POLYGON  4.0150 1.2500 3.0850 1.2500 3.0850 1.8700 2.9650 1.8700 2.9650 0.8600 2.9050 0.8600
                 2.9050 0.7400 3.1450 0.7400 3.1450 0.8600 3.0850 0.8600 3.0850 1.1300 4.0150 1.1300 ;
        POLYGON  2.6450 1.8700 2.5250 1.8700 2.5250 1.8600 0.9200 1.8600 0.9200 1.7700 0.4350 1.7700
                 0.4350 1.6500 0.9200 1.6500 0.9200 0.9600 0.8050 0.9600 0.8050 0.6800 0.9250 0.6800
                 0.9250 0.8400 1.0400 0.8400 1.0400 1.7400 2.3650 1.7400 2.3650 0.8000 2.4250 0.8000
                 2.4250 0.6800 2.5450 0.6800 2.5450 0.9200 2.4850 0.9200 2.4850 1.6300 2.6450 1.6300 ;
        POLYGON  1.9850 1.1600 1.8650 1.1600 1.8650 0.9000 1.3450 0.9000 1.3450 1.5000 1.4650 1.5000
                 1.4650 1.6200 1.2250 1.6200 1.2250 0.6600 1.1950 0.6600 1.1950 0.4200 1.3150 0.4200
                 1.3150 0.5400 1.3450 0.5400 1.3450 0.7800 1.9850 0.7800 ;
    END
END DFFTRX4

MACRO DFFTRX2
    CLASS CORE ;
    FOREIGN DFFTRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2950 0.8850 0.4150 1.3700 ;
        RECT  0.0700 0.8850 0.4150 1.3400 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.0700 1.0900 1.4350 ;
        RECT  0.8350 0.9150 0.9550 1.2900 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7900 1.0050 6.0300 1.1800 ;
        RECT  5.8700 0.8000 6.0200 1.1800 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6100 1.3600 6.7300 2.0100 ;
        RECT  6.5700 0.7400 6.6900 1.4800 ;
        RECT  6.4500 0.7400 6.6900 1.1450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.4100 0.7400 7.6500 0.8600 ;
        RECT  7.4500 1.3000 7.5700 2.0100 ;
        RECT  7.4100 0.7400 7.5300 1.4200 ;
        RECT  7.3200 0.8850 7.5300 1.1450 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.9500 -0.1800 8.0700 0.3800 ;
        RECT  6.9300 -0.1800 7.1700 0.3800 ;
        RECT  5.9700 -0.1800 6.2100 0.3800 ;
        RECT  4.7400 -0.1800 4.8600 0.7600 ;
        RECT  2.9600 0.3500 3.2000 0.4700 ;
        RECT  2.9600 -0.1800 3.0800 0.4700 ;
        RECT  0.9100 -0.1800 1.0300 0.7500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.8700 1.3600 7.9900 2.7900 ;
        RECT  7.0300 1.3600 7.1500 2.7900 ;
        RECT  6.1900 1.3600 6.3100 2.7900 ;
        RECT  4.7800 2.1600 5.0200 2.2800 ;
        RECT  4.7800 2.1600 4.9000 2.7900 ;
        RECT  2.9800 2.2300 3.2200 2.7900 ;
        RECT  1.0350 2.0100 1.1550 2.7900 ;
        RECT  0.1350 1.4900 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.5500 1.1800 8.4700 1.1800 8.4700 1.6000 8.3500 1.6000 8.3500 1.1800 7.6700 1.1800
                 7.6700 1.0600 8.4300 1.0600 8.4300 0.6800 8.5500 0.6800 ;
        POLYGON  8.4500 0.5200 8.3100 0.5200 8.3100 0.6200 6.9850 0.6200 6.9850 1.2400 6.8650 1.2400
                 6.8650 0.6200 6.3300 0.6200 6.3300 1.2400 6.2100 1.2400 6.2100 0.6200 5.2800 0.6200
                 5.2800 0.7600 5.3000 0.7600 5.3000 1.6800 5.5000 1.6800 5.5000 1.8000 5.1800 1.8000
                 5.1800 1.5200 4.8200 1.5200 4.8200 1.2800 4.9400 1.2800 4.9400 1.4000 5.1800 1.4000
                 5.1800 0.8800 5.1600 0.8800 5.1600 0.5000 8.1900 0.5000 8.1900 0.4000 8.4500 0.4000 ;
        POLYGON  5.8300 2.0400 4.5150 2.0400 4.5150 2.1100 4.1050 2.1100 4.1050 2.2500 3.8650 2.2500
                 3.8650 2.1100 2.6600 2.1100 2.6600 2.2500 2.4200 2.2500 2.4200 2.1300 2.5400 2.1300
                 2.5400 1.9900 4.3950 1.9900 4.3950 1.9200 5.7100 1.9200 5.7100 1.4800 5.5500 1.4800
                 5.5500 0.8600 5.4900 0.8600 5.4900 0.7400 5.7300 0.7400 5.7300 0.8600 5.6700 0.8600
                 5.6700 1.3600 5.8300 1.3600 ;
        POLYGON  5.0600 1.1200 4.7000 1.1200 4.7000 1.7300 4.2600 1.7300 4.2600 1.8700 4.1400 1.8700
                 4.1400 1.6100 4.5800 1.6100 4.5800 1.1200 4.0400 1.1200 4.0400 0.6200 4.1600 0.6200
                 4.1600 1.0000 5.0600 1.0000 ;
        POLYGON  4.4600 1.4900 3.8000 1.4900 3.8000 1.3100 3.7200 1.3100 3.7200 1.0700 3.8000 1.0700
                 3.8000 0.5000 3.4400 0.5000 3.4400 0.7100 2.7200 0.7100 2.7200 0.5000 2.1100 0.5000
                 2.1100 1.3700 2.2000 1.3700 2.2000 1.4900 1.9600 1.4900 1.9600 1.3700 1.9900 1.3700
                 1.9900 0.5000 1.5800 0.5000 1.5800 0.5100 1.4500 0.5100 1.4500 1.3700 1.6000 1.3700
                 1.6000 1.6100 1.4800 1.6100 1.4800 1.4900 1.3300 1.4900 1.3300 0.3900 1.4600 0.3900
                 1.4600 0.3800 2.4000 0.3800 2.4000 0.3600 2.6400 0.3600 2.6400 0.3800 2.8400 0.3800
                 2.8400 0.5900 3.3200 0.5900 3.3200 0.3800 3.9200 0.3800 3.9200 1.3700 4.4600 1.3700 ;
        POLYGON  3.6800 0.9500 3.6000 0.9500 3.6000 1.6300 3.6400 1.6300 3.6400 1.8700 3.5200 1.8700
                 3.5200 1.7500 3.4800 1.7500 3.4800 1.4900 2.7800 1.4900 2.7800 1.3700 3.4800 1.3700
                 3.4800 0.8300 3.5600 0.8300 3.5600 0.6200 3.6800 0.6200 ;
        POLYGON  3.3600 1.2500 2.4600 1.2500 2.4600 1.8700 2.3400 1.8700 2.3400 0.8000 2.2600 0.8000
                 2.2600 0.6800 2.5000 0.6800 2.5000 0.8000 2.4600 0.8000 2.4600 1.1300 3.3600 1.1300 ;
        POLYGON  2.0400 1.8700 1.9200 1.8700 1.9200 1.8500 0.5550 1.8500 0.5550 1.6100 0.5350 1.6100
                 0.5350 0.7650 0.2700 0.7650 0.2700 0.5100 0.3900 0.5100 0.3900 0.6450 0.6550 0.6450
                 0.6550 1.4900 0.6750 1.4900 0.6750 1.7300 1.7200 1.7300 1.7200 0.6200 1.8400 0.6200
                 1.8400 1.6300 2.0400 1.6300 ;
    END
END DFFTRX2

MACRO DFFTRX1
    CLASS CORE ;
    FOREIGN DFFTRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8400 1.3400 2.1400 1.4600 ;
        RECT  2.0200 1.2200 2.1400 1.4600 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.8400 1.3400 1.9600 1.7250 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0800 1.0900 7.2000 1.3300 ;
        RECT  6.7400 1.1750 7.2000 1.2950 ;
        RECT  6.7400 1.1750 6.8900 1.4350 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.4100 1.0100 7.5600 1.2500 ;
        RECT  7.3200 0.8850 7.4950 1.1450 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3800 1.3000 1.5000 2.2100 ;
        RECT  1.3800 0.6200 1.5000 0.8600 ;
        RECT  1.3600 0.7400 1.4800 1.4200 ;
        RECT  1.2300 0.8850 1.4800 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  6.9600 -0.1800 7.0800 0.9100 ;
        RECT  4.8300 -0.1800 5.0700 0.3200 ;
        RECT  3.2300 -0.1800 3.3500 0.9000 ;
        RECT  1.8000 -0.1800 1.9200 0.7300 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.8000 1.8100 7.9200 2.7900 ;
        RECT  6.9000 2.2300 7.0200 2.7900 ;
        RECT  4.8300 2.1600 5.0700 2.2800 ;
        RECT  4.8300 2.1600 4.9500 2.7900 ;
        RECT  3.1100 2.1600 3.3500 2.2800 ;
        RECT  3.1100 2.1600 3.2300 2.7900 ;
        RECT  1.8000 1.8450 1.9200 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.8000 1.4900 7.5000 1.4900 7.5000 2.1100 6.0550 2.1100 6.0550 1.9800 6.0300 1.9800
                 6.0300 1.5100 6.1900 1.5100 6.1900 0.9000 6.1300 0.9000 6.1300 0.6600 6.2500 0.6600
                 6.2500 0.7800 6.3100 0.7800 6.3100 1.6300 6.1500 1.6300 6.1500 1.8600 6.1750 1.8600
                 6.1750 1.9900 7.3800 1.9900 7.3800 1.3700 7.6800 1.3700 7.6800 0.6700 7.8000 0.6700 ;
        POLYGON  6.6600 0.9100 6.6200 0.9100 6.6200 1.8700 6.3600 1.8700 6.3600 1.7500 6.5000 1.7500
                 6.5000 0.7900 6.5400 0.7900 6.5400 0.6700 6.4300 0.6700 6.4300 0.5400 6.0100 0.5400
                 6.0100 1.2700 6.0700 1.2700 6.0700 1.3900 5.8300 1.3900 5.8300 1.2700 5.8900 1.2700
                 5.8900 0.5400 5.3100 0.5400 5.3100 0.5600 4.2300 0.5600 4.2300 1.0000 4.3700 1.0000
                 4.3700 1.2400 4.2300 1.2400 4.2300 1.4000 3.8300 1.4000 3.8300 1.5200 3.7100 1.5200
                 3.7100 1.2800 4.1100 1.2800 4.1100 0.4400 5.1900 0.4400 5.1900 0.4200 5.3700 0.4200
                 5.3700 0.3800 5.6100 0.3800 5.6100 0.4200 6.5500 0.4200 6.5500 0.5500 6.6600 0.5500 ;
        POLYGON  5.7700 0.8400 5.7100 0.8400 5.7100 1.6200 5.7300 1.6200 5.7300 1.8600 5.6100 1.8600
                 5.6100 1.7400 5.5900 1.7400 5.5900 1.4800 4.7300 1.4800 4.7300 1.3600 5.5900 1.3600
                 5.5900 0.8400 5.5300 0.8400 5.5300 0.7200 5.7700 0.7200 ;
        POLYGON  5.6300 2.2400 5.1950 2.2400 5.1950 2.0400 4.2550 2.0400 4.2550 2.2400 4.0150 2.2400
                 4.0150 2.0400 2.2800 2.0400 2.2800 0.6800 2.4000 0.6800 2.4000 1.9200 5.3150 1.9200
                 5.3150 2.1200 5.6300 2.1200 ;
        POLYGON  5.2700 1.1600 4.6100 1.1600 4.6100 1.8000 4.3500 1.8000 4.3500 1.6800 4.4900 1.6800
                 4.4900 0.8400 4.3500 0.8400 4.3500 0.7200 4.6100 0.7200 4.6100 1.0400 5.2700 1.0400 ;
        POLYGON  4.0500 1.8000 3.8100 1.8000 3.8100 1.7600 3.4700 1.7600 3.4700 1.4000 2.9500 1.4000
                 2.9500 1.5200 2.8300 1.5200 2.8300 1.2800 3.4700 1.2800 3.4700 1.0400 3.8700 1.0400
                 3.8700 0.6600 3.9900 0.6600 3.9900 1.1600 3.5900 1.1600 3.5900 1.6400 3.9300 1.6400
                 3.9300 1.6800 4.0500 1.6800 ;
        POLYGON  3.3500 1.1600 2.7100 1.1600 2.7100 1.6800 2.8700 1.6800 2.8700 1.8000 2.5900 1.8000
                 2.5900 0.7800 2.6700 0.7800 2.6700 0.6600 2.5700 0.6600 2.5700 0.5600 2.1600 0.5600
                 2.1600 1.1000 1.8400 1.1000 1.8400 1.1800 1.6000 1.1800 1.6000 0.9800 2.0400 0.9800
                 2.0400 0.4400 2.6900 0.4400 2.6900 0.5400 2.7900 0.5400 2.7900 0.9000 2.7100 0.9000
                 2.7100 1.0400 3.3500 1.0400 ;
        POLYGON  1.1100 1.0800 1.0950 1.0800 1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000
                 0.3750 1.0800 0.9750 1.0800 0.9750 0.9600 0.9900 0.9600 0.9900 0.6800 1.1100 0.6800 ;
    END
END DFFTRX1

MACRO DFFSXL
    CLASS CORE ;
    FOREIGN DFFSXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1350 1.2200 3.4650 1.4350 ;
        RECT  3.0150 1.2200 3.4650 1.4100 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0350 1.2200 8.1550 1.5100 ;
        RECT  7.9000 1.1750 8.0500 1.4750 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4800 1.0400 8.6300 1.4350 ;
        RECT  8.4800 0.8350 8.6000 1.4350 ;
        END
    END CK
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6600 1.4850 1.5800 ;
        RECT  1.2300 0.8850 1.4850 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.3750 -0.1800 8.4950 0.3800 ;
        RECT  6.6050 -0.1800 6.8450 0.3200 ;
        RECT  3.2950 -0.1800 3.4150 0.4000 ;
        RECT  1.8450 -0.1800 1.9650 0.3800 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.1950 1.6800 8.3150 2.7900 ;
        RECT  6.9550 2.2000 7.0750 2.7900 ;
        RECT  4.3750 2.2900 4.6150 2.7900 ;
        RECT  3.4750 2.0500 3.5950 2.7900 ;
        RECT  2.5150 1.7300 2.6350 2.7900 ;
        RECT  1.8450 1.9800 1.9650 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.8700 1.6750 8.7350 1.6750 8.7350 1.8000 8.6150 1.8000 8.6150 1.5550 8.7500 1.5550
                 8.7500 0.9000 8.7350 0.9000 8.7350 0.6600 8.1350 0.6600 8.1350 0.5400 7.5150 0.5400
                 7.5150 1.4600 7.3950 1.4600 7.3950 0.5600 5.6750 0.5600 5.6750 1.4600 5.5550 1.4600
                 5.5550 0.5600 5.1950 0.5600 5.1950 0.5200 5.0750 0.5200 5.0750 0.4000 5.3150 0.4000
                 5.3150 0.4400 6.2450 0.4400 6.2450 0.4000 6.4850 0.4000 6.4850 0.4400 7.3950 0.4400
                 7.3950 0.4200 7.7550 0.4200 7.7550 0.4000 7.9950 0.4000 7.9950 0.4200 8.2550 0.4200
                 8.2550 0.5400 8.8550 0.5400 8.8550 0.7800 8.8700 0.7800 ;
        POLYGON  7.7550 1.7000 7.6750 1.7000 7.6750 1.9400 6.8350 1.9400 6.8350 2.2200 4.7350 2.2200
                 4.7350 2.1700 4.0550 2.1700 4.0550 2.0500 4.8550 2.0500 4.8550 2.1000 6.7150 2.1000
                 6.7150 1.8200 7.5550 1.8200 7.5550 1.5800 7.6350 1.5800 7.6350 0.6600 7.7550 0.6600 ;
        POLYGON  7.1950 1.4600 7.0750 1.4600 7.0750 1.1800 6.2450 1.1800 6.2450 1.6200 6.3550 1.6200
                 6.3550 1.7400 6.1150 1.7400 6.1150 1.6200 6.1250 1.6200 6.1250 1.2600 6.0350 1.2600
                 6.0350 1.0200 6.1250 1.0200 6.1250 0.7200 6.3650 0.7200 6.3650 0.8400 6.2450 0.8400
                 6.2450 1.0600 7.1950 1.0600 ;
        POLYGON  6.9150 1.4200 6.7950 1.4200 6.7950 1.7000 6.5950 1.7000 6.5950 1.9800 5.7850 1.9800
                 5.7850 1.9600 5.0650 1.9600 5.0650 1.6000 4.8000 1.6000 4.8000 1.5700 4.1350 1.5700
                 4.1350 1.6900 3.8950 1.6900 3.8950 1.5700 4.0150 1.5700 4.0150 1.4500 4.2750 1.4500
                 4.2750 0.6800 4.3950 0.6800 4.3950 1.4500 4.9200 1.4500 4.9200 1.4800 5.1850 1.4800
                 5.1850 1.8400 5.7850 1.8400 5.7850 1.5800 5.7950 1.5800 5.7950 0.6800 5.9150 0.6800
                 5.9150 1.7000 5.9050 1.7000 5.9050 1.8600 6.4750 1.8600 6.4750 1.5800 6.6750 1.5800
                 6.6750 1.3000 6.9150 1.3000 ;
        POLYGON  5.5450 1.7200 5.3050 1.7200 5.3050 1.1600 4.5150 1.1600 4.5150 0.5600 4.1550 0.5600
                 4.1550 0.7200 4.0350 0.7200 4.0350 1.1000 2.1850 1.1000 2.1850 1.2200 2.0650 1.2200
                 2.0650 0.9800 3.9150 0.9800 3.9150 0.6000 4.0350 0.6000 4.0350 0.4400 4.6350 0.4400
                 4.6350 1.0400 5.3050 1.0400 5.3050 0.8600 5.1950 0.8600 5.1950 0.7400 5.4350 0.7400
                 5.4350 0.8600 5.4250 0.8600 5.4250 1.6000 5.5450 1.6000 ;
        POLYGON  4.9550 0.9200 4.8350 0.9200 4.8350 0.7200 4.7550 0.7200 4.7550 0.3600 4.8750 0.3600
                 4.8750 0.6000 4.9550 0.6000 ;
        POLYGON  4.9450 1.8400 4.8250 1.8400 4.8250 1.9300 2.9950 1.9300 2.9950 1.6300 3.1150 1.6300
                 3.1150 1.8100 4.7050 1.8100 4.7050 1.7200 4.9450 1.7200 ;
        POLYGON  3.9150 0.4800 3.7950 0.4800 3.7950 0.7400 2.7750 0.7400 2.7750 0.8600 2.5350 0.8600
                 2.5350 0.7400 2.6550 0.7400 2.6550 0.6200 3.6750 0.6200 3.6750 0.3600 3.9150 0.3600 ;
        POLYGON  2.8950 1.3700 2.4250 1.3700 2.4250 1.4600 2.3250 1.4600 2.3250 1.5800 2.2050 1.5800
                 2.2050 1.4600 1.8250 1.4600 1.8250 1.2000 1.6050 1.2000 1.6050 1.0800 1.8250 1.0800
                 1.8250 0.7200 2.3850 0.7200 2.3850 0.8400 1.9450 0.8400 1.9450 1.3400 2.3050 1.3400
                 2.3050 1.2500 2.8950 1.2500 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFSXL

MACRO DFFSX4
    CLASS CORE ;
    FOREIGN DFFSX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4100 1.0000 0.5300 1.4850 ;
        RECT  0.3600 1.0000 0.5300 1.4550 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7500 1.0000 0.8700 1.3800 ;
        RECT  0.6500 1.1300 0.8000 1.5000 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.4500 1.2550 5.5700 1.4950 ;
        RECT  4.7100 1.2550 5.5700 1.3750 ;
        RECT  4.7700 0.3950 4.8900 1.3750 ;
        RECT  4.7100 1.1750 4.8600 1.4350 ;
        RECT  3.3850 0.3950 4.8900 0.5150 ;
        RECT  2.9050 0.9800 3.5050 1.1000 ;
        RECT  3.3850 0.3950 3.5050 1.1000 ;
        RECT  2.9050 0.3600 3.0250 1.1000 ;
        RECT  2.7850 0.3600 3.0250 0.4800 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.9700 1.4400 8.0900 2.2100 ;
        RECT  6.8900 0.8000 7.9700 0.9200 ;
        RECT  7.8500 0.6800 7.9700 0.9200 ;
        RECT  7.7900 1.4400 8.0900 1.5600 ;
        RECT  7.3100 1.3200 7.9100 1.4400 ;
        RECT  7.3100 1.1750 7.4700 1.4400 ;
        RECT  7.1300 1.4400 7.4300 1.5600 ;
        RECT  7.3100 0.8000 7.4300 1.5600 ;
        RECT  7.1300 1.4400 7.2500 2.2100 ;
        RECT  6.8900 0.6800 7.0100 0.9200 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8100 0.8000 9.8900 0.9200 ;
        RECT  9.7700 0.6800 9.8900 0.9200 ;
        RECT  9.6500 1.4400 9.7700 2.2100 ;
        RECT  9.4700 1.4400 9.7700 1.5600 ;
        RECT  8.8000 1.3200 9.5900 1.4400 ;
        RECT  8.8100 0.6800 8.9300 2.2100 ;
        RECT  8.7700 1.1750 8.9300 1.4350 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.2500 -0.1800 10.3700 0.7300 ;
        RECT  9.2300 -0.1800 9.4700 0.3200 ;
        RECT  8.2700 -0.1800 8.5100 0.3200 ;
        RECT  7.3100 -0.1800 7.5500 0.3200 ;
        RECT  6.4100 -0.1800 6.5300 0.8200 ;
        RECT  5.5700 -0.1800 5.6900 0.8750 ;
        RECT  3.1450 -0.1800 3.2650 0.8600 ;
        RECT  1.9950 -0.1800 2.2350 0.3200 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.0700 1.6000 10.1900 2.7900 ;
        RECT  9.2300 1.5600 9.3500 2.7900 ;
        RECT  8.3900 1.5600 8.5100 2.7900 ;
        RECT  7.5500 1.5600 7.6700 2.7900 ;
        RECT  6.7100 1.5600 6.8300 2.7900 ;
        RECT  5.7500 1.9400 5.9900 2.1500 ;
        RECT  5.7500 1.9400 5.8700 2.7900 ;
        RECT  4.8500 2.1800 5.0900 2.3000 ;
        RECT  4.8500 2.1800 4.9700 2.7900 ;
        RECT  2.8300 2.2800 3.0700 2.7900 ;
        RECT  1.9300 2.1000 2.0500 2.7900 ;
        RECT  0.5900 1.6200 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.7900 1.4800 10.6100 1.4800 10.6100 2.2100 10.4900 2.2100 10.4900 1.4800
                 9.9150 1.4800 9.9150 1.2400 10.0350 1.2400 10.0350 1.3600 10.6700 1.3600
                 10.6700 0.6800 10.7900 0.6800 ;
        POLYGON  10.3950 1.2400 10.2750 1.2400 10.2750 0.9700 10.0100 0.9700 10.0100 0.5600
                 6.7700 0.5600 6.7700 1.0400 6.9700 1.0400 6.9700 1.2800 6.8500 1.2800 6.8500 1.1600
                 6.3500 1.1600 6.3500 2.2100 6.2300 2.2100 6.2300 1.1350 5.0100 1.1350 5.0100 1.0150
                 5.9900 1.0150 5.9900 0.6800 6.1100 0.6800 6.1100 0.9400 6.6500 0.9400 6.6500 0.4400
                 10.1300 0.4400 10.1300 0.8500 10.3950 0.8500 ;
        POLYGON  6.0900 1.5900 5.8100 1.5900 5.8100 1.8200 4.2200 1.8200 4.2200 2.0900 4.1000 2.0900
                 4.1000 1.7000 4.4700 1.7000 4.4700 0.9350 4.5300 0.9350 4.5300 0.6350 4.6500 0.6350
                 4.6500 1.0550 4.5900 1.0550 4.5900 1.7000 5.6900 1.7000 5.6900 1.4700 5.9700 1.4700
                 5.9700 1.3500 6.0900 1.3500 ;
        RECT  4.4600 1.9400 5.5700 2.0600 ;
        POLYGON  4.3500 1.5800 3.8000 1.5800 3.8000 2.1300 3.6800 2.1300 3.6800 1.9200 3.0700 1.9200
                 3.0700 1.7400 2.4100 1.7400 2.4100 1.5000 2.4250 1.5000 2.4250 1.0200 1.7750 1.0200
                 1.7750 0.9000 2.3050 0.9000 2.3050 0.6800 2.4250 0.6800 2.4250 0.8400 2.5450 0.8400
                 2.5450 1.6200 3.1900 1.6200 3.1900 1.8000 3.6800 1.8000 3.6800 1.4600 4.2300 1.4600
                 4.2300 0.8150 4.0500 0.8150 4.0500 0.6950 4.3500 0.6950 ;
        POLYGON  4.1100 1.3400 3.5500 1.3400 3.5500 1.6800 3.3100 1.6800 3.3100 1.5600 3.4300 1.5600
                 3.4300 1.3400 2.6650 1.3400 2.6650 0.7200 2.5450 0.7200 2.5450 0.5600 1.6350 0.5600
                 1.6350 0.9800 1.5150 0.9800 1.5150 0.4400 2.6650 0.4400 2.6650 0.6000 2.7850 0.6000
                 2.7850 1.2200 3.6250 1.2200 3.6250 0.6800 3.7450 0.6800 3.7450 1.2200 3.9900 1.2200
                 3.9900 0.9600 4.1100 0.9600 ;
        POLYGON  3.3900 2.1600 2.8300 2.1600 2.8300 1.9800 1.5100 1.9800 1.5100 2.2000 1.3900 2.2000
                 1.3900 1.9800 0.9900 1.9800 0.9900 0.8800 0.2400 0.8800 0.2400 1.5750 0.2900 1.5750
                 0.2900 1.8150 0.1700 1.8150 0.1700 1.6950 0.1200 1.6950 0.1200 0.6400 0.1350 0.6400
                 0.1350 0.4000 0.2550 0.4000 0.2550 0.7600 1.0350 0.7600 1.0350 0.7400 1.1550 0.7400
                 1.1550 0.9800 1.1100 0.9800 1.1100 1.8600 2.9500 1.8600 2.9500 2.0400 3.3900 2.0400 ;
        POLYGON  2.3050 1.3600 1.3950 1.3600 1.3950 1.6200 1.3500 1.6200 1.3500 1.7400 1.2300 1.7400
                 1.2300 1.5000 1.2750 1.5000 1.2750 0.4000 1.3950 0.4000 1.3950 1.2400 2.3050 1.2400 ;
    END
END DFFSX4

MACRO DFFSX2
    CLASS CORE ;
    FOREIGN DFFSX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0500 0.5100 1.5200 ;
        RECT  0.3900 1.0200 0.5100 1.5200 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0800 0.8350 1.5100 ;
        RECT  0.6500 1.1450 0.8000 1.5600 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5800 1.4650 5.7300 1.7250 ;
        RECT  5.5800 1.1300 5.7000 1.7250 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6100 1.1750 7.7600 1.4350 ;
        RECT  7.6350 1.1750 7.7550 2.1600 ;
        RECT  7.6100 0.7400 7.7300 1.4350 ;
        RECT  7.4550 0.7400 7.7300 0.8600 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4150 0.7400 8.6550 0.8600 ;
        RECT  8.4800 1.1750 8.6300 1.4350 ;
        RECT  8.4800 0.7400 8.6000 1.4350 ;
        RECT  8.4750 1.2950 8.5950 2.1600 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.8950 -0.1800 9.1350 0.3200 ;
        RECT  7.9350 -0.1800 8.1750 0.3800 ;
        RECT  6.9750 -0.1800 7.2150 0.3800 ;
        RECT  5.4050 0.4100 5.6450 0.5300 ;
        RECT  5.5250 -0.1800 5.6450 0.5300 ;
        RECT  1.6150 -0.1800 1.8550 0.3200 ;
        RECT  0.6150 -0.1800 0.7350 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.8950 1.5100 9.0150 2.7900 ;
        RECT  8.0550 1.5100 8.1750 2.7900 ;
        RECT  7.2150 1.6400 7.3350 2.7900 ;
        RECT  6.4050 2.0900 6.5250 2.7900 ;
        RECT  5.6650 2.0900 5.7850 2.7900 ;
        RECT  4.6400 2.2900 4.8800 2.7900 ;
        RECT  1.9550 2.2000 2.0750 2.7900 ;
        RECT  0.6550 1.6800 0.7750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.4950 0.8600 9.4350 0.8600 9.4350 1.7500 9.3150 1.7500 9.3150 1.2900 8.7500 1.2900
                 8.7500 1.1700 9.3150 1.1700 9.3150 0.8600 9.2550 0.8600 9.2550 0.7400 9.4950 0.7400 ;
        POLYGON  9.4150 0.6200 8.0000 0.6200 8.0000 1.2400 7.8800 1.2400 7.8800 0.6200 7.3350 0.6200
                 7.3350 1.0600 7.4550 1.0600 7.4550 1.1800 7.1150 1.1800 7.1150 1.5200 6.9750 1.5200
                 6.9750 2.1000 6.7350 2.1000 6.7350 1.7000 6.8550 1.7000 6.8550 1.4000 6.9950 1.4000
                 6.9950 1.0400 6.1550 1.0400 6.1550 0.9200 6.5550 0.9200 6.5550 0.6800 6.6750 0.6800
                 6.6750 0.9200 7.2150 0.9200 7.2150 0.5000 9.2950 0.5000 9.2950 0.3600 9.4150 0.3600 ;
        POLYGON  6.8750 1.2800 5.9150 1.2800 5.9150 1.0100 5.4600 1.0100 5.4600 1.2400 4.6250 1.2400
                 4.6250 1.1200 5.3400 1.1200 5.3400 0.8900 6.0350 0.8900 6.0350 1.1600 6.8750 1.1600 ;
        POLYGON  6.3450 0.7200 6.2250 0.7200 6.2250 0.7700 5.0650 0.7700 5.0650 0.4800 4.5850 0.4800
                 4.5850 0.6000 4.2650 0.6000 4.2650 0.8200 4.0250 0.8200 4.0250 0.7000 4.1450 0.7000
                 4.1450 0.4800 4.4650 0.4800 4.4650 0.3600 5.1850 0.3600 5.1850 0.6500 6.1050 0.6500
                 6.1050 0.6000 6.3450 0.6000 ;
        POLYGON  6.1450 1.9650 5.3400 1.9650 5.3400 1.9300 4.2650 1.9300 4.2650 1.8200 4.1450 1.8200
                 4.1450 1.7000 4.3850 1.7000 4.3850 1.8100 5.4600 1.8100 5.4600 1.8450 6.0250 1.8450
                 6.0250 1.5700 6.1450 1.5700 ;
        POLYGON  5.3050 1.6900 5.1850 1.6900 5.1850 1.5700 4.5050 1.5700 4.5050 1.5800 4.0250 1.5800
                 4.0250 1.9800 2.4350 1.9800 2.4350 1.4000 2.1950 1.4000 2.1950 1.2800 2.5550 1.2800
                 2.5550 1.8600 3.1650 1.8600 3.1650 1.7400 3.1250 1.7400 3.1250 0.7600 3.1850 0.7600
                 3.1850 0.6400 3.3050 0.6400 3.3050 0.8800 3.2450 0.8800 3.2450 1.6200 3.2850 1.6200
                 3.2850 1.8600 3.9050 1.8600 3.9050 1.4600 4.3850 1.4600 4.3850 0.7200 4.7050 0.7200
                 4.7050 0.6000 4.9450 0.6000 4.9450 0.7200 4.8250 0.7200 4.8250 0.8400 4.5050 0.8400
                 4.5050 1.4500 5.3050 1.4500 ;
        POLYGON  5.2200 2.1700 4.3050 2.1700 4.3050 2.2200 2.1950 2.2200 2.1950 2.0400 1.4150 2.0400
                 1.4150 1.8000 1.3350 1.8000 1.3350 0.8400 1.2150 0.8400 1.2150 0.7200 1.4550 0.7200
                 1.4550 1.6800 1.5350 1.6800 1.5350 1.9200 2.3150 1.9200 2.3150 2.1000 4.1850 2.1000
                 4.1850 2.0500 5.2200 2.0500 ;
        POLYGON  4.2650 1.3400 3.7850 1.3400 3.7850 1.7000 3.5250 1.7000 3.5250 1.5800 3.6650 1.5800
                 3.6650 0.6400 3.7850 0.6400 3.7850 1.2200 4.2650 1.2200 ;
        POLYGON  4.0050 0.4800 3.8850 0.4800 3.8850 0.5000 3.5450 0.5000 3.5450 1.1200 3.4850 1.1200
                 3.4850 1.4400 3.3650 1.4400 3.3650 1.0000 3.4250 1.0000 3.4250 0.5000 2.2200 0.5000
                 2.2200 0.6000 1.6950 0.6000 1.6950 1.4600 1.5750 1.4600 1.5750 0.6000 1.0950 0.6000
                 1.0950 1.0000 1.1550 1.0000 1.1550 1.2400 0.9750 1.2400 0.9750 0.9000 0.2400 0.9000
                 0.2400 1.6400 0.3550 1.6400 0.3550 1.8800 0.2350 1.8800 0.2350 1.7600 0.1200 1.7600
                 0.1200 0.7800 0.1350 0.7800 0.1350 0.6600 0.2550 0.6600 0.2550 0.7800 0.9750 0.7800
                 0.9750 0.4800 2.1000 0.4800 2.1000 0.3800 3.7650 0.3800 3.7650 0.3600 4.0050 0.3600 ;
        POLYGON  3.0050 1.2200 2.8550 1.2200 2.8550 1.6200 2.9150 1.6200 2.9150 1.7400 2.6750 1.7400
                 2.6750 1.6200 2.7350 1.6200 2.7350 1.1600 2.0750 1.1600 2.0750 1.1800 1.8350 1.1800
                 1.8350 1.0400 2.7350 1.0400 2.7350 0.7200 2.9750 0.7200 2.9750 0.8400 2.8550 0.8400
                 2.8550 0.9800 3.0050 0.9800 ;
    END
END DFFSX2

MACRO DFFSX1
    CLASS CORE ;
    FOREIGN DFFSX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1350 1.2000 3.4650 1.4150 ;
        RECT  3.0150 1.2000 3.4650 1.3900 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0350 1.2200 8.1550 1.5100 ;
        RECT  7.9000 1.1750 8.0500 1.4750 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.4800 1.0400 8.6300 1.4350 ;
        RECT  8.4950 0.8350 8.6150 1.4350 ;
        END
    END CK
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6600 1.4850 1.9900 ;
        RECT  1.2300 0.8850 1.4850 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.3750 -0.1800 8.4950 0.3800 ;
        RECT  6.6050 -0.1800 6.8450 0.3200 ;
        RECT  3.2950 -0.1800 3.4150 0.3800 ;
        RECT  1.8450 -0.1800 1.9650 0.3800 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.1950 1.6800 8.3150 2.7900 ;
        RECT  6.9550 2.2000 7.0750 2.7900 ;
        RECT  4.3750 2.2900 4.6150 2.7900 ;
        RECT  3.4750 2.0500 3.5950 2.7900 ;
        RECT  2.5150 1.7300 2.6350 2.7900 ;
        RECT  1.7850 1.3400 1.9050 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.8700 1.6750 8.7350 1.6750 8.7350 1.8000 8.6150 1.8000 8.6150 1.5550 8.7500 1.5550
                 8.7500 0.9000 8.7350 0.9000 8.7350 0.6600 8.1350 0.6600 8.1350 0.5400 7.5150 0.5400
                 7.5150 1.4600 7.3950 1.4600 7.3950 0.5600 5.6750 0.5600 5.6750 1.4600 5.5550 1.4600
                 5.5550 0.5600 5.1950 0.5600 5.1950 0.5200 5.0750 0.5200 5.0750 0.4000 5.3150 0.4000
                 5.3150 0.4400 6.2450 0.4400 6.2450 0.4000 6.4850 0.4000 6.4850 0.4400 7.3950 0.4400
                 7.3950 0.4200 7.7550 0.4200 7.7550 0.4000 7.9950 0.4000 7.9950 0.4200 8.2550 0.4200
                 8.2550 0.5400 8.8550 0.5400 8.8550 0.7800 8.8700 0.7800 ;
        POLYGON  7.7550 1.7000 7.6750 1.7000 7.6750 1.9400 6.8350 1.9400 6.8350 2.2200 4.7350 2.2200
                 4.7350 2.1700 4.0550 2.1700 4.0550 2.0500 4.8550 2.0500 4.8550 2.1000 6.7150 2.1000
                 6.7150 1.8200 7.5550 1.8200 7.5550 1.5800 7.6350 1.5800 7.6350 0.6600 7.7550 0.6600 ;
        POLYGON  7.1950 1.4600 7.0750 1.4600 7.0750 1.1800 6.2450 1.1800 6.2450 1.6200 6.3550 1.6200
                 6.3550 1.7400 6.1150 1.7400 6.1150 1.6200 6.1250 1.6200 6.1250 1.2600 6.0350 1.2600
                 6.0350 1.0200 6.1250 1.0200 6.1250 0.7200 6.3650 0.7200 6.3650 0.8400 6.2450 0.8400
                 6.2450 1.0600 7.1950 1.0600 ;
        POLYGON  6.9150 1.4200 6.7950 1.4200 6.7950 1.7000 6.5950 1.7000 6.5950 1.9800 5.7850 1.9800
                 5.7850 1.9600 5.0650 1.9600 5.0650 1.6000 4.8000 1.6000 4.8000 1.5700 4.1350 1.5700
                 4.1350 1.6900 3.8950 1.6900 3.8950 1.5700 4.0150 1.5700 4.0150 1.4500 4.2750 1.4500
                 4.2750 0.6600 4.3950 0.6600 4.3950 1.4500 4.9200 1.4500 4.9200 1.4800 5.1850 1.4800
                 5.1850 1.8400 5.7850 1.8400 5.7850 1.5800 5.7950 1.5800 5.7950 0.6800 5.9150 0.6800
                 5.9150 1.7000 5.9050 1.7000 5.9050 1.8600 6.4750 1.8600 6.4750 1.5800 6.6750 1.5800
                 6.6750 1.3000 6.9150 1.3000 ;
        POLYGON  5.5450 1.7200 5.3050 1.7200 5.3050 1.1600 4.5150 1.1600 4.5150 0.5400 4.1550 0.5400
                 4.1550 0.7200 4.0350 0.7200 4.0350 1.0800 2.3850 1.0800 2.3850 1.2200 2.2650 1.2200
                 2.2650 0.9600 3.9150 0.9600 3.9150 0.6000 4.0350 0.6000 4.0350 0.4200 4.6350 0.4200
                 4.6350 1.0400 5.3050 1.0400 5.3050 0.8600 5.1950 0.8600 5.1950 0.7400 5.4350 0.7400
                 5.4350 0.8600 5.4250 0.8600 5.4250 1.6000 5.5450 1.6000 ;
        POLYGON  4.9550 0.9200 4.8350 0.9200 4.8350 0.6000 4.7550 0.6000 4.7550 0.3600 4.8750 0.3600
                 4.8750 0.4800 4.9550 0.4800 ;
        POLYGON  4.9450 1.8400 4.8250 1.8400 4.8250 1.9300 2.9950 1.9300 2.9950 1.6300 3.1150 1.6300
                 3.1150 1.8100 4.7050 1.8100 4.7050 1.7200 4.9450 1.7200 ;
        POLYGON  3.9150 0.4800 3.7950 0.4800 3.7950 0.7200 2.7750 0.7200 2.7750 0.8400 2.5350 0.8400
                 2.5350 0.7200 2.6550 0.7200 2.6550 0.6000 3.6750 0.6000 3.6750 0.3600 3.9150 0.3600 ;
        POLYGON  2.8950 1.3700 2.6250 1.3700 2.6250 1.4600 2.3250 1.4600 2.3250 1.5800 2.2050 1.5800
                 2.2050 1.4600 2.0250 1.4600 2.0250 1.2000 1.6050 1.2000 1.6050 1.0800 2.0250 1.0800
                 2.0250 0.7200 2.3850 0.7200 2.3850 0.8400 2.1450 0.8400 2.1450 1.3400 2.5050 1.3400
                 2.5050 1.2500 2.8950 1.2500 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFSX1

MACRO DFFSRXL
    CLASS CORE ;
    FOREIGN DFFSRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8750 1.4800 2.1150 1.6400 ;
        RECT  1.7550 1.5200 2.0150 1.7150 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5900 1.2300 7.6500 1.3500 ;
        RECT  6.0500 1.1200 6.7100 1.2400 ;
        RECT  6.0500 0.4000 6.1700 1.2400 ;
        RECT  5.0850 0.4000 6.1700 0.5200 ;
        RECT  3.2800 1.1600 5.2050 1.2800 ;
        RECT  5.0850 0.4000 5.2050 1.2800 ;
        RECT  4.9450 0.9400 5.2050 1.2800 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3500 1.1200 9.5550 1.4350 ;
        RECT  9.3500 1.0700 9.5250 1.4350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5100 1.0400 10.6600 1.4500 ;
        RECT  10.5250 1.0400 10.6450 1.5250 ;
        END
    END CK
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 0.6800 1.4850 0.9200 ;
        RECT  1.3550 1.3200 1.4750 2.0900 ;
        RECT  1.3350 0.8000 1.4550 1.4400 ;
        RECT  1.2300 0.8850 1.4550 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.7050 -0.1800 10.8250 0.9200 ;
        RECT  9.4500 -0.1800 9.5700 0.8900 ;
        RECT  7.7500 -0.1800 7.9900 0.3200 ;
        RECT  3.0750 -0.1800 3.1950 0.7800 ;
        RECT  1.7850 -0.1800 1.9050 0.9200 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.7650 1.5700 10.8850 2.7900 ;
        RECT  9.5900 2.1700 9.7100 2.7900 ;
        RECT  8.0500 2.2900 8.2900 2.7900 ;
        RECT  6.5700 2.2900 6.8100 2.7900 ;
        RECT  4.2600 1.8800 4.3800 2.7900 ;
        RECT  2.8800 2.2800 3.1200 2.7900 ;
        RECT  1.7750 1.9700 1.8950 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.4050 0.9200 10.3900 0.9200 10.3900 1.5700 10.4050 1.5700 10.4050 2.0350
                 10.1100 2.0350 10.1100 2.1300 9.8700 2.1300 9.8700 2.0500 9.4700 2.0500 9.4700 2.1700
                 6.4650 2.1700 6.4650 2.1200 5.5500 2.1200 5.5500 2.0000 6.5850 2.0000 6.5850 2.0500
                 9.3500 2.0500 9.3500 1.9300 9.8700 1.9300 9.8700 1.9150 10.2850 1.9150 10.2850 1.6900
                 10.2700 1.6900 10.2700 0.8000 10.2850 0.8000 10.2850 0.6800 10.4050 0.6800 ;
        POLYGON  10.0150 1.7950 9.8950 1.7950 9.8950 1.6750 9.2300 1.6750 9.2300 1.9300 6.7800 1.9300
                 6.7800 1.8800 5.4300 1.8800 5.4300 2.0800 4.8700 2.0800 4.8700 1.9600 5.3100 1.9600
                 5.3100 1.7600 5.5650 1.7600 5.5650 1.0800 5.5700 1.0800 5.5700 0.9600 5.6900 0.9600
                 5.6900 1.2000 5.6850 1.2000 5.6850 1.7600 6.9000 1.7600 6.9000 1.8100 8.3700 1.8100
                 8.3700 0.9700 8.4900 0.9700 8.4900 1.8100 9.1100 1.8100 9.1100 1.4500 8.9500 1.4500
                 8.9500 1.1900 9.0700 1.1900 9.0700 1.3300 9.2300 1.3300 9.2300 1.5550 9.8700 1.5550
                 9.8700 0.6500 9.9900 0.6500 9.9900 1.5550 10.0150 1.5550 ;
        POLYGON  8.9900 1.6900 8.6100 1.6900 8.6100 0.6500 7.6300 0.6500 7.6300 0.6000 7.3100 0.6000
                 7.3100 0.5200 7.1900 0.5200 7.1900 0.4000 7.4300 0.4000 7.4300 0.4800 7.7500 0.4800
                 7.7500 0.5300 8.7300 0.5300 8.7300 1.5700 8.9900 1.5700 ;
        POLYGON  8.1500 1.2300 8.0300 1.2300 8.0300 1.1100 7.8900 1.1100 7.8900 1.5900 7.5100 1.5900
                 7.5100 1.6900 7.2700 1.6900 7.2700 1.5900 6.0450 1.5900 6.0450 1.6400 5.8050 1.6400
                 5.8050 1.5200 5.8100 1.5200 5.8100 0.6400 5.9300 0.6400 5.9300 1.4700 7.7700 1.4700
                 7.7700 1.1100 6.8300 1.1100 6.8300 1.0000 6.7100 1.0000 6.7100 0.6600 6.8300 0.6600
                 6.8300 0.8800 6.9500 0.8800 6.9500 0.9900 8.1500 0.9900 ;
        POLYGON  7.5100 0.8400 7.0700 0.8400 7.0700 0.7600 6.9500 0.7600 6.9500 0.5400 6.4100 0.5400
                 6.4100 0.9000 6.2900 0.9000 6.2900 0.4200 7.0700 0.4200 7.0700 0.6400 7.1900 0.6400
                 7.1900 0.7200 7.5100 0.7200 ;
        POLYGON  5.4500 0.8800 5.4450 0.8800 5.4450 1.5800 5.1900 1.5800 5.1900 1.7000 5.0700 1.7000
                 5.0700 1.5200 2.9200 1.5200 2.9200 1.2600 3.0400 1.2600 3.0400 1.4000 5.3250 1.4000
                 5.3250 0.7600 5.3300 0.7600 5.3300 0.6400 5.4500 0.6400 ;
        POLYGON  4.9650 0.8200 4.7550 0.8200 4.7550 0.9600 4.0350 0.9600 4.0350 0.7200 3.8550 0.7200
                 3.8550 0.6000 4.1550 0.6000 4.1550 0.8400 4.6350 0.8400 4.6350 0.7000 4.9650 0.7000 ;
        POLYGON  4.8300 1.7600 4.1300 1.7600 4.1300 1.8100 3.3600 1.8100 3.3600 1.6900 4.0100 1.6900
                 4.0100 1.6400 4.8300 1.6400 ;
        POLYGON  4.5150 0.7200 4.2750 0.7200 4.2750 0.4800 3.7350 0.4800 3.7350 0.5400 3.6150 0.5400
                 3.6150 0.7800 3.4950 0.7800 3.4950 0.4200 3.6150 0.4200 3.6150 0.3600 4.3950 0.3600
                 4.3950 0.6000 4.5150 0.6000 ;
        POLYGON  4.1000 2.2500 3.3300 2.2500 3.3300 2.1600 2.3150 2.1600 2.3150 2.2100 2.1950 2.2100
                 2.1950 1.9700 2.2650 1.9700 2.2650 0.6800 2.3850 0.6800 2.3850 2.0400 3.4500 2.0400
                 3.4500 2.1300 4.1000 2.1300 ;
        POLYGON  3.8800 1.0400 2.7750 1.0400 2.7750 1.7000 2.6250 1.7000 2.6250 1.8200 2.5050 1.8200
                 2.5050 1.5800 2.6550 1.5800 2.6550 0.5600 2.1450 0.5600 2.1450 1.2000 1.5750 1.2000
                 1.5750 1.0800 2.0250 1.0800 2.0250 0.4400 2.7750 0.4400 2.7750 0.9200 3.8800 0.9200 ;
        POLYGON  1.2150 1.5800 1.0950 1.5800 1.0950 1.4600 0.9750 1.4600 0.9750 1.2000 0.3750 1.2000
                 0.3750 1.0800 0.9750 1.0800 0.9750 0.6800 1.0950 0.6800 1.0950 1.3400 1.2150 1.3400 ;
    END
END DFFSRXL

MACRO DFFSRX4
    CLASS CORE ;
    FOREIGN DFFSRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.2100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 1.0650 0.5100 1.5500 ;
        RECT  0.3600 1.0650 0.5100 1.5200 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0250 1.4100 1.2650 1.5550 ;
        RECT  0.8850 1.5000 1.1450 1.6700 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6750 1.1200 4.9550 1.2400 ;
        RECT  4.6550 1.2300 4.9500 1.3800 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2000 1.2300 5.4950 1.3800 ;
        RECT  5.2150 1.1200 5.4950 1.3800 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.9150 0.7400 11.1150 0.8600 ;
        RECT  10.9350 1.4200 11.0550 2.1900 ;
        RECT  10.6350 1.4200 11.0550 1.5400 ;
        RECT  9.9300 1.3000 10.7550 1.4200 ;
        RECT  9.9750 0.7400 10.0950 2.1900 ;
        RECT  9.9300 1.1750 10.0950 1.4350 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.8350 0.7400 13.0350 0.8600 ;
        RECT  12.6550 1.4200 12.7750 2.1900 ;
        RECT  12.4750 1.4200 12.7750 1.5400 ;
        RECT  11.9900 1.3000 12.5950 1.4200 ;
        RECT  11.8150 1.4200 12.1100 1.5400 ;
        RECT  11.9900 0.7400 12.1100 1.5400 ;
        RECT  11.9600 0.7400 12.1100 1.1450 ;
        RECT  11.8150 1.4200 11.9350 2.1900 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.2100 0.1800 ;
        RECT  13.3950 -0.1800 13.5150 0.7300 ;
        RECT  12.3150 -0.1800 12.5550 0.3800 ;
        RECT  11.3550 -0.1800 11.5950 0.3800 ;
        RECT  10.3950 -0.1800 10.6350 0.3800 ;
        RECT  9.3150 0.6400 9.5550 0.7600 ;
        RECT  9.3150 -0.1800 9.4350 0.7600 ;
        RECT  8.5350 -0.1800 8.6550 0.8600 ;
        RECT  5.0350 0.6400 5.2750 0.7600 ;
        RECT  5.1550 -0.1800 5.2750 0.7600 ;
        RECT  2.3850 -0.1800 2.6250 0.3600 ;
        RECT  0.6250 -0.1800 0.7450 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.2100 2.7900 ;
        RECT  13.0750 1.5400 13.1950 2.7900 ;
        RECT  12.2350 1.5400 12.3550 2.7900 ;
        RECT  11.3950 1.5400 11.5150 2.7900 ;
        RECT  10.3950 1.5400 10.5150 2.7900 ;
        RECT  9.5550 1.6000 9.6750 2.7900 ;
        RECT  8.7100 1.7600 8.8300 2.7900 ;
        RECT  7.6500 1.8800 7.7700 2.7900 ;
        RECT  4.8950 1.9800 5.0150 2.7900 ;
        RECT  4.7750 1.9800 5.0150 2.1000 ;
        RECT  3.2150 2.1600 3.3350 2.7900 ;
        RECT  3.0950 2.1600 3.3350 2.2800 ;
        RECT  2.2450 2.1600 2.4850 2.2800 ;
        RECT  2.2450 2.1600 2.3650 2.7900 ;
        RECT  0.9650 1.7900 1.0850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.9350 0.9200 13.7750 0.9200 13.7750 1.4200 13.6150 1.4200 13.6150 2.1900
                 13.4950 2.1900 13.4950 1.4200 12.8950 1.4200 12.8950 1.2800 13.1350 1.2800
                 13.1350 1.3000 13.6550 1.3000 13.6550 0.8000 13.8150 0.8000 13.8150 0.6800
                 13.9350 0.6800 ;
        POLYGON  13.5350 1.1800 13.2950 1.1800 13.2950 0.9700 13.1550 0.9700 13.1550 0.6200
                 9.7950 0.6200 9.7950 1.0000 9.2300 1.0000 9.2300 1.2800 9.8100 1.2800 9.8100 1.4000
                 9.2500 1.4000 9.2500 2.1200 9.1300 2.1200 9.1300 1.4000 9.1100 1.4000 9.1100 1.1400
                 7.9950 1.1400 7.9950 1.0200 8.9550 1.0200 8.9550 0.6800 9.0750 0.6800 9.0750 0.8800
                 9.6750 0.8800 9.6750 0.5000 13.2750 0.5000 13.2750 0.8500 13.4150 0.8500
                 13.4150 1.0600 13.5350 1.0600 ;
        POLYGON  8.9900 1.5200 6.5250 1.5200 6.5250 1.8900 6.4050 1.8900 6.4050 0.9200 6.3850 0.9200
                 6.3850 0.6800 6.5050 0.6800 6.5050 0.8000 6.5250 0.8000 6.5250 1.4000 8.8700 1.4000
                 8.8700 1.2600 8.9900 1.2600 ;
        POLYGON  8.4700 1.9400 8.2050 1.9400 8.2050 1.7600 7.5300 1.7600 7.5300 1.8100 6.7650 1.8100
                 6.7650 1.6900 7.4100 1.6900 7.4100 1.6400 8.3250 1.6400 8.3250 1.8200 8.4700 1.8200 ;
        POLYGON  8.2350 0.8600 8.1150 0.8600 8.1150 0.5000 7.5750 0.5000 7.5750 0.6800 7.4550 0.6800
                 7.4550 0.8000 7.2150 0.8000 7.2150 0.6800 7.3350 0.6800 7.3350 0.5600 7.4550 0.5600
                 7.4550 0.3800 8.2350 0.3800 ;
        POLYGON  7.8150 1.0400 6.9750 1.0400 6.9750 0.9200 6.8850 0.9200 6.8850 0.6800 7.0050 0.6800
                 7.0050 0.8000 7.0950 0.8000 7.0950 0.9200 7.6950 0.9200 7.6950 0.6200 7.8150 0.6200 ;
        POLYGON  7.6150 1.2800 6.7350 1.2800 6.7350 1.1600 6.6450 1.1600 6.6450 0.5600 5.7050 0.5600
                 5.7050 0.7400 5.7350 0.7400 5.7350 1.6200 5.6150 1.6200 5.6150 1.0000 4.7950 1.0000
                 4.7950 0.5000 4.3800 0.5000 4.3800 0.4800 3.9950 0.4800 3.9950 0.3600 4.5000 0.3600
                 4.5000 0.3800 4.9150 0.3800 4.9150 0.8800 5.5750 0.8800 5.5750 0.6200 5.5850 0.6200
                 5.5850 0.4400 6.7650 0.4400 6.7650 1.0400 6.8550 1.0400 6.8550 1.1600 7.6150 1.1600 ;
        POLYGON  6.7850 2.2500 5.6650 2.2500 5.6650 2.1300 5.1350 2.1300 5.1350 1.8600 4.0550 1.8600
                 4.0550 1.5600 2.7250 1.5600 2.7250 1.4400 2.8450 1.4400 2.8450 0.9400 2.0050 0.9400
                 2.0050 1.2200 1.8850 1.2200 1.8850 0.8200 2.8450 0.8200 2.8450 0.7200 3.1050 0.7200
                 3.1050 0.8400 2.9650 0.8400 2.9650 1.4400 4.1750 1.4400 4.1750 1.7400 5.2550 1.7400
                 5.2550 2.0100 5.7850 2.0100 5.7850 2.1300 6.1650 2.1300 6.1650 1.2800 6.1250 1.2800
                 6.1250 1.0400 6.2850 1.0400 6.2850 2.1300 6.7850 2.1300 ;
        POLYGON  6.0850 0.9200 6.0050 0.9200 6.0050 1.7700 6.0450 1.7700 6.0450 2.0100 5.9250 2.0100
                 5.9250 1.8900 5.3750 1.8900 5.3750 1.6200 4.2950 1.6200 4.2950 1.5000 4.4150 1.5000
                 4.4150 1.3200 3.2750 1.3200 3.2750 0.5000 3.0600 0.5000 3.0600 0.6000 2.1450 0.6000
                 2.1450 0.5200 2.0250 0.5200 2.0250 0.4000 2.2650 0.4000 2.2650 0.4800 2.9400 0.4800
                 2.9400 0.3800 3.8750 0.3800 3.8750 0.6800 4.3150 0.6800 4.3150 0.8000 3.7550 0.8000
                 3.7550 0.5000 3.3950 0.5000 3.3950 1.2000 4.5350 1.2000 4.5350 1.5000 5.4950 1.5000
                 5.4950 1.7700 5.8850 1.7700 5.8850 0.8000 5.9650 0.8000 5.9650 0.6800 6.0850 0.6800 ;
        POLYGON  4.6750 1.0000 4.5550 1.0000 4.5550 1.0400 3.5150 1.0400 3.5150 0.6200 3.6350 0.6200
                 3.6350 0.9200 4.4350 0.9200 4.4350 0.8800 4.5550 0.8800 4.5550 0.6200 4.6750 0.6200 ;
        POLYGON  4.6550 2.2500 4.0800 2.2500 4.0800 2.1000 3.8150 2.1000 3.8150 1.8000 2.4850 1.8000
                 2.4850 1.4800 1.6450 1.4800 1.6450 0.5400 1.2850 0.5400 1.2850 1.2400 1.1650 1.2400
                 1.1650 0.9450 0.2400 0.9450 0.2400 1.6700 0.5850 1.6700 0.5850 1.9100 0.4650 1.9100
                 0.4650 1.7900 0.1200 1.7900 0.1200 0.7800 0.1450 0.7800 0.1450 0.6600 0.2650 0.6600
                 0.2650 0.8250 1.1650 0.8250 1.1650 0.4200 1.7650 0.4200 1.7650 1.3600 2.4850 1.3600
                 2.4850 1.0600 2.6250 1.0600 2.6250 1.3000 2.6050 1.3000 2.6050 1.6800 3.9350 1.6800
                 3.9350 1.9800 4.2000 1.9800 4.2000 2.1300 4.6550 2.1300 ;
        POLYGON  3.6950 2.1600 3.4550 2.1600 3.4550 2.0400 1.6050 2.0400 1.6050 1.8000 1.4050 1.8000
                 1.4050 0.6600 1.5250 0.6600 1.5250 1.6800 1.7250 1.6800 1.7250 1.9200 3.5750 1.9200
                 3.5750 2.0400 3.6950 2.0400 ;
    END
END DFFSRX4

MACRO DFFSRX2
    CLASS CORE ;
    FOREIGN DFFSRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.0500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2850 1.0200 0.4050 1.2600 ;
        RECT  0.0700 1.0200 0.4050 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2600 1.5350 1.4500 ;
        RECT  1.1750 1.2300 1.4350 1.4500 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.8976  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 7.4800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 1.2000 3.1750 1.4700 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1650 1.1200 10.4250 1.3800 ;
        RECT  10.1750 1.0200 10.4150 1.3800 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.9150 0.6800 11.0350 2.0300 ;
        RECT  10.8000 1.4650 11.0350 1.7250 ;
        RECT  10.8300 1.3800 11.0350 1.7250 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.7150 0.7400 12.0550 0.8600 ;
        RECT  11.7550 1.3200 11.8750 2.0300 ;
        RECT  11.6700 1.1750 11.8350 1.4350 ;
        RECT  11.7150 0.7400 11.8350 1.4400 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.0500 0.1800 ;
        RECT  12.2950 -0.1800 12.5350 0.3200 ;
        RECT  11.3350 -0.1800 11.5750 0.3200 ;
        RECT  10.3750 -0.1800 10.6150 0.3200 ;
        RECT  9.2650 -0.1800 9.3850 0.8300 ;
        RECT  2.5950 0.7200 2.8350 0.8400 ;
        RECT  2.5950 -0.1800 2.7150 0.8400 ;
        RECT  1.4350 -0.1800 1.5550 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.0500 2.7900 ;
        RECT  12.1750 1.3800 12.2950 2.7900 ;
        RECT  11.3350 1.3800 11.4550 2.7900 ;
        RECT  10.4950 1.5000 10.6150 2.7900 ;
        RECT  9.1850 2.1300 9.3050 2.7900 ;
        RECT  9.0650 2.1300 9.3050 2.2500 ;
        RECT  6.3850 1.8800 6.6250 2.0000 ;
        RECT  6.3850 1.8800 6.5050 2.7900 ;
        RECT  4.1650 2.0000 4.4050 2.1200 ;
        RECT  4.1650 2.0000 4.2850 2.7900 ;
        RECT  2.9050 2.1300 3.0250 2.7900 ;
        RECT  1.1950 1.8700 1.3150 2.7900 ;
        RECT  0.1350 1.9800 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  12.9750 0.8600 12.8550 0.8600 12.8550 1.2000 12.7150 1.2000 12.7150 1.6200
                 12.5950 1.6200 12.5950 1.2000 11.9550 1.2000 11.9550 1.0800 12.7350 1.0800
                 12.7350 0.7400 12.9750 0.7400 ;
        POLYGON  12.8950 0.5200 12.7750 0.5200 12.7750 0.5600 11.2750 0.5600 11.2750 1.2600
                 11.1550 1.2600 11.1550 0.5600 10.7750 0.5600 10.7750 1.2600 10.6550 1.2600
                 10.6550 0.6000 9.8050 0.6000 9.8050 1.5900 9.7850 1.5900 9.7850 2.0100 9.6650 2.0100
                 9.6650 1.4700 9.6850 1.4700 9.6850 1.1100 8.6250 1.1100 8.6250 0.9900 9.6850 0.9900
                 9.6850 0.4800 10.6550 0.4800 10.6550 0.4400 12.6550 0.4400 12.6550 0.4000
                 12.8950 0.4000 ;
        POLYGON  10.2550 0.8400 10.0450 0.8400 10.0450 1.6200 10.1950 1.6200 10.1950 2.2500
                 9.4250 2.2500 9.4250 2.0100 6.9850 2.0100 6.9850 1.5200 6.1650 1.5200 6.1650 1.4000
                 7.1050 1.4000 7.1050 1.8900 9.5450 1.8900 9.5450 2.1300 10.0750 2.1300 10.0750 1.7400
                 9.9250 1.7400 9.9250 0.7200 10.2550 0.7200 ;
        POLYGON  9.5650 1.3500 7.4650 1.3500 7.4650 1.0400 5.6450 1.0400 5.6450 1.6400 5.6050 1.6400
                 5.6050 1.7600 5.4850 1.7600 5.4850 1.5200 5.5250 1.5200 5.5250 0.6200 5.6450 0.6200
                 5.6450 0.9200 7.5850 0.9200 7.5850 1.2300 9.5650 1.2300 ;
        POLYGON  9.0250 0.7700 8.7250 0.7700 8.7250 0.5300 8.1850 0.5300 8.1850 0.7700 7.9450 0.7700
                 7.9450 0.6500 8.0650 0.6500 8.0650 0.4100 8.8450 0.4100 8.8450 0.6500 9.0250 0.6500 ;
        POLYGON  8.9450 2.2500 6.7450 2.2500 6.7450 1.7600 6.2650 1.7600 6.2650 2.0000 5.7050 2.0000
                 5.7050 2.2400 4.5250 2.2400 4.5250 1.8800 4.0450 1.8800 4.0450 2.2500 3.1650 2.2500
                 3.1650 2.1300 3.9250 2.1300 3.9250 1.7600 4.6450 1.7600 4.6450 2.1200 5.5850 2.1200
                 5.5850 1.8800 6.1450 1.8800 6.1450 1.6400 6.8650 1.6400 6.8650 2.1300 8.9450 2.1300 ;
        POLYGON  8.8250 1.7700 7.2250 1.7700 7.2250 1.2800 6.0250 1.2800 6.0250 1.7600 5.9050 1.7600
                 5.9050 1.1600 7.3450 1.1600 7.3450 1.6500 8.8250 1.6500 ;
        POLYGON  8.6050 0.7700 8.4250 0.7700 8.4250 1.0100 7.7050 1.0100 7.7050 0.8000 5.8850 0.8000
                 5.8850 0.6800 7.8250 0.6800 7.8250 0.8900 8.3050 0.8900 8.3050 0.6500 8.6050 0.6500 ;
        POLYGON  5.8450 0.4800 5.4050 0.4800 5.4050 1.3000 5.3650 1.3000 5.3650 2.0000 4.7650 2.0000
                 4.7650 1.6400 3.8050 1.6400 3.8050 2.0100 2.5850 2.0100 2.5850 2.2300 2.4950 2.2300
                 2.4950 2.2500 2.2550 2.2500 2.2550 2.2300 1.9350 2.2300 1.9350 1.2300 1.7750 1.2300
                 1.7750 1.1100 1.0550 1.1100 1.0550 0.9900 1.1950 0.9900 1.1950 0.4900 0.6850 0.4900
                 0.6850 0.8000 0.6950 0.8000 0.6950 1.5800 0.5750 1.5800 0.5750 0.9200 0.5650 0.9200
                 0.5650 0.3700 1.3150 0.3700 1.3150 0.9900 1.8950 0.9900 1.8950 1.0400 2.0550 1.0400
                 2.0550 2.1100 2.4650 2.1100 2.4650 1.8900 3.6850 1.8900 3.6850 1.5200 4.8850 1.5200
                 4.8850 1.8800 5.2450 1.8800 5.2450 1.1800 5.2850 1.1800 5.2850 0.3600 5.8450 0.3600 ;
        POLYGON  5.1650 1.0600 5.1250 1.0600 5.1250 1.7600 5.0050 1.7600 5.0050 1.4000 3.4450 1.4000
                 3.4450 1.6500 3.5650 1.6500 3.5650 1.7700 3.3250 1.7700 3.3250 1.7100 2.6550 1.7100
                 2.6550 1.2900 2.7750 1.2900 2.7750 1.5900 3.3250 1.5900 3.3250 1.2800 3.6550 1.2800
                 3.6550 0.9200 3.6050 0.9200 3.6050 0.6600 3.7250 0.6600 3.7250 0.8000 3.7750 0.8000
                 3.7750 1.2800 5.0050 1.2800 5.0050 0.9400 5.0450 0.9400 5.0450 0.6200 5.1650 0.6200 ;
        POLYGON  4.1450 0.9000 4.0250 0.9000 4.0250 0.5400 3.4850 0.5400 3.4850 0.7200 3.3650 0.7200
                 3.3650 0.8400 3.1250 0.8400 3.1250 0.7200 3.2450 0.7200 3.2450 0.6000 3.3650 0.6000
                 3.3650 0.4200 4.1450 0.4200 ;
        POLYGON  3.5350 1.1600 3.2950 1.1600 3.2950 1.0800 2.2950 1.0800 2.2950 1.9900 2.1750 1.9900
                 2.1750 0.9200 2.0150 0.9200 2.0150 0.6600 2.1350 0.6600 2.1350 0.8000 2.2950 0.8000
                 2.2950 0.9600 3.4150 0.9600 3.4150 1.0400 3.5350 1.0400 ;
        POLYGON  1.8150 1.6900 0.9350 1.6900 0.9350 1.8200 0.8950 1.8200 0.8950 2.0900 0.7750 2.0900
                 0.7750 1.7000 0.8150 1.7000 0.8150 0.7300 0.9550 0.7300 0.9550 0.6100 1.0750 0.6100
                 1.0750 0.8500 0.9350 0.8500 0.9350 1.5700 1.6950 1.5700 1.6950 1.4100 1.8150 1.4100 ;
    END
END DFFSRX2

MACRO DFFSRX1
    CLASS CORE ;
    FOREIGN DFFSRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.7300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9150 1.1000 2.1550 1.2250 ;
        RECT  1.7550 1.2250 2.0350 1.3800 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5850 1.2400 7.6450 1.3600 ;
        RECT  6.0450 1.1200 6.7050 1.2400 ;
        RECT  6.0450 0.4000 6.1650 1.2400 ;
        RECT  5.0850 0.4000 6.1650 0.5200 ;
        RECT  3.3150 1.2400 5.2050 1.3600 ;
        RECT  5.0850 0.4000 5.2050 1.3600 ;
        RECT  4.9450 0.9400 5.2050 1.0900 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3500 1.1750 9.5000 1.4350 ;
        RECT  9.1850 1.1200 9.4700 1.2400 ;
        RECT  9.1850 1.0000 9.3050 1.2400 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.3350 1.0150 10.6600 1.1500 ;
        RECT  10.5100 0.8850 10.6600 1.1500 ;
        RECT  10.3350 1.0150 10.4550 1.2600 ;
        END
    END CK
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2744  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3750 0.5000 1.4950 0.7400 ;
        RECT  1.3650 1.5850 1.4850 2.0300 ;
        RECT  1.2300 1.4650 1.4350 1.7250 ;
        RECT  1.3150 0.6200 1.4350 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.7300 0.1800 ;
        RECT  10.4750 -0.1800 10.5950 0.4000 ;
        RECT  9.1850 -0.1800 9.3050 0.8800 ;
        RECT  7.7450 -0.1800 7.9850 0.3200 ;
        RECT  3.0550 0.6600 3.2950 0.7800 ;
        RECT  3.1750 -0.1800 3.2950 0.7800 ;
        RECT  1.7950 -0.1800 1.9150 0.7400 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.7300 2.7900 ;
        RECT  10.4750 1.9700 10.5950 2.7900 ;
        RECT  9.4250 2.1000 9.5450 2.7900 ;
        RECT  7.7450 2.2900 7.9850 2.7900 ;
        RECT  6.4250 2.2000 6.6650 2.7900 ;
        RECT  4.3750 2.0500 4.4950 2.7900 ;
        RECT  2.9950 1.9600 3.1150 2.7900 ;
        RECT  1.7850 1.5000 1.9050 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.2150 1.9700 10.1750 1.9700 10.1750 2.0900 10.0550 2.0900 10.0550 1.9800
                 9.3050 1.9800 9.3050 2.1800 8.1050 2.1800 8.1050 2.1700 6.7850 2.1700 6.7850 2.0800
                 5.5450 2.0800 5.5450 1.9600 6.9050 1.9600 6.9050 2.0500 8.2250 2.0500 8.2250 2.0600
                 9.1850 2.0600 9.1850 1.8600 9.6550 1.8600 9.6550 1.8400 9.8950 1.8400 9.8950 1.8600
                 10.0550 1.8600 10.0550 1.8500 10.0950 1.8500 10.0950 0.9200 10.0550 0.9200
                 10.0550 0.6800 10.1750 0.6800 10.1750 0.8000 10.2150 0.8000 ;
        POLYGON  9.9750 1.7000 9.8550 1.7000 9.8550 1.6750 9.0650 1.6750 9.0650 1.9400 8.3450 1.9400
                 8.3450 1.9300 7.0250 1.9300 7.0250 1.8400 5.4250 1.8400 5.4250 2.1600 4.8650 2.1600
                 4.8650 2.0400 5.3050 2.0400 5.3050 1.7200 5.5650 1.7200 5.5650 0.9600 5.6850 0.9600
                 5.6850 1.7200 7.1450 1.7200 7.1450 1.8100 8.2450 1.8100 8.2450 0.9800 8.3650 0.9800
                 8.3650 1.8100 8.4650 1.8100 8.4650 1.8200 8.9450 1.8200 8.9450 1.4400 8.8250 1.4400
                 8.8250 1.2000 9.0650 1.2000 9.0650 1.5550 9.6650 1.5550 9.6650 0.6600 9.7850 0.6600
                 9.7850 1.4600 9.9750 1.4600 ;
        POLYGON  8.8250 1.7000 8.5850 1.7000 8.5850 0.9000 8.4850 0.9000 8.4850 0.6600 7.6250 0.6600
                 7.6250 0.5600 7.3050 0.5600 7.3050 0.5200 7.1850 0.5200 7.1850 0.4000 7.4250 0.4000
                 7.4250 0.4400 7.7450 0.4400 7.7450 0.5400 8.6050 0.5400 8.6050 0.7800 8.7050 0.7800
                 8.7050 1.5800 8.8250 1.5800 ;
        POLYGON  8.0250 1.2400 7.8850 1.2400 7.8850 1.6000 7.5050 1.6000 7.5050 1.6900 7.2650 1.6900
                 7.2650 1.6000 5.8050 1.6000 5.8050 0.6400 5.9250 0.6400 5.9250 1.4800 7.7650 1.4800
                 7.7650 1.1200 6.8250 1.1200 6.8250 1.0000 6.7050 1.0000 6.7050 0.6600 6.8250 0.6600
                 6.8250 0.8800 6.9450 0.8800 6.9450 1.0000 8.0250 1.0000 ;
        POLYGON  7.5050 0.8400 7.0650 0.8400 7.0650 0.7600 6.9450 0.7600 6.9450 0.5400 6.4050 0.5400
                 6.4050 0.9000 6.2850 0.9000 6.2850 0.4200 7.0650 0.4200 7.0650 0.6400 7.1850 0.6400
                 7.1850 0.7200 7.5050 0.7200 ;
        POLYGON  5.4450 1.6000 5.1850 1.6000 5.1850 1.7800 5.0650 1.7800 5.0650 1.6000 2.9750 1.6000
                 2.9750 1.3600 3.0950 1.3600 3.0950 1.4800 5.3250 1.4800 5.3250 0.6400 5.4450 0.6400 ;
        POLYGON  4.9650 0.8200 4.8250 0.8200 4.8250 1.0800 3.9950 1.0800 3.9950 0.8400 3.9550 0.8400
                 3.9550 0.6000 4.0750 0.6000 4.0750 0.7200 4.1150 0.7200 4.1150 0.9600 4.7050 0.9600
                 4.7050 0.7000 4.9650 0.7000 ;
        POLYGON  4.8250 1.8400 4.7050 1.8400 4.7050 1.9300 3.4750 1.9300 3.4750 1.8100 4.5850 1.8100
                 4.5850 1.7200 4.8250 1.7200 ;
        POLYGON  4.4950 0.8400 4.3750 0.8400 4.3750 0.7200 4.2350 0.7200 4.2350 0.4800 3.8250 0.4800
                 3.8250 0.6000 3.6550 0.6000 3.6550 0.8400 3.5350 0.8400 3.5350 0.4800 3.7050 0.4800
                 3.7050 0.3600 4.3550 0.3600 4.3550 0.6000 4.4950 0.6000 ;
        POLYGON  4.2150 2.2500 3.9750 2.2500 3.9750 2.1700 3.2350 2.1700 3.2350 1.8400 2.8750 1.8400
                 2.8750 2.2500 2.2050 2.2500 2.2050 1.3800 2.2750 1.3800 2.2750 0.6000 2.3950 0.6000
                 2.3950 1.5000 2.3250 1.5000 2.3250 2.1300 2.7550 2.1300 2.7550 1.7200 3.3550 1.7200
                 3.3550 2.0500 4.0950 2.0500 4.0950 2.1300 4.2150 2.1300 ;
        POLYGON  3.8750 1.1200 2.8150 1.1200 2.8150 1.6000 2.6350 1.6000 2.6350 2.0100 2.5150 2.0100
                 2.5150 1.4800 2.6950 1.4800 2.6950 0.4800 2.1550 0.4800 2.1550 0.9800 1.7950 0.9800
                 1.7950 1.1050 1.5550 1.1050 1.5550 0.8600 2.0350 0.8600 2.0350 0.3600 2.8150 0.3600
                 2.8150 1.0000 3.8750 1.0000 ;
        POLYGON  1.1100 1.5800 0.9900 1.5800 0.9900 1.4600 0.9850 1.4600 0.9850 1.1800 0.3750 1.1800
                 0.3750 1.0600 0.9850 1.0600 0.9850 0.6800 1.1050 0.6800 1.1050 1.3400 1.1100 1.3400 ;
    END
END DFFSRX1

MACRO DFFSRHQX8
    CLASS CORE ;
    FOREIGN DFFSRHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.6300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 1.4650 2.7750 2.2100 ;
        RECT  2.6550 0.6800 2.7750 1.0050 ;
        RECT  2.6350 0.8850 2.7550 1.5850 ;
        RECT  0.0700 1.0050 2.7550 1.1250 ;
        RECT  1.8150 0.6800 1.9350 2.2100 ;
        RECT  0.9750 0.6800 1.0950 2.2050 ;
        RECT  0.1350 0.6800 0.2550 2.2050 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 1.0200 5.1500 1.4350 ;
        RECT  5.0000 0.9200 5.1200 1.4350 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3200 2.1300 9.8250 2.2500 ;
        RECT  9.3200 1.7600 9.4400 2.2500 ;
        RECT  8.5650 1.7600 9.4400 1.8800 ;
        RECT  7.0850 2.1300 8.6850 2.2500 ;
        RECT  8.5650 1.7600 8.6850 2.2500 ;
        RECT  7.0850 1.7600 7.2050 2.2500 ;
        RECT  6.2350 1.7600 7.2050 1.8800 ;
        RECT  5.7050 1.8900 6.3550 2.0100 ;
        RECT  6.2350 1.7600 6.3550 2.0100 ;
        RECT  5.7050 1.2300 5.8250 2.0100 ;
        RECT  5.5800 1.1750 5.7300 1.4350 ;
        RECT  5.6100 1.1100 5.7300 1.4350 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.9050 0.8950 12.1650 1.1300 ;
        RECT  11.8250 1.0100 12.0650 1.2200 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.1200 1.1600 13.2700 1.5800 ;
        RECT  13.1250 1.0400 13.2450 1.5800 ;
        END
    END CK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.6300 0.1800 ;
        RECT  13.3750 -0.1800 13.4950 0.4000 ;
        RECT  12.0450 -0.1800 12.2850 0.3200 ;
        RECT  10.5050 -0.1800 10.6250 0.6800 ;
        RECT  5.2050 -0.1800 5.4450 0.3200 ;
        RECT  3.9150 -0.1800 4.0350 0.6900 ;
        RECT  3.0750 -0.1800 3.1950 0.6900 ;
        RECT  2.2350 -0.1800 2.3550 0.6700 ;
        RECT  1.3950 -0.1800 1.5150 0.6700 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.6300 2.7900 ;
        RECT  13.3000 1.7000 13.4200 2.7900 ;
        RECT  12.0250 1.5800 12.1450 2.7900 ;
        RECT  10.5200 1.8600 10.6400 2.7900 ;
        RECT  10.4000 1.8600 10.6400 2.0000 ;
        RECT  8.9250 2.0000 9.0450 2.7900 ;
        RECT  8.8050 2.0000 9.0450 2.1200 ;
        RECT  6.7250 2.0000 6.9650 2.1200 ;
        RECT  6.7250 2.0000 6.8450 2.7900 ;
        RECT  5.2250 1.7950 5.3450 2.7900 ;
        RECT  5.1050 1.7950 5.3450 1.9150 ;
        RECT  3.9150 1.5600 4.0350 2.7900 ;
        RECT  3.0750 1.5600 3.1950 2.7900 ;
        RECT  2.2350 1.4650 2.3550 2.7900 ;
        RECT  1.3950 1.4650 1.5150 2.7900 ;
        RECT  0.5550 1.4650 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.0950 0.9200 13.0050 0.9200 13.0050 1.0400 13.0000 1.0400 13.0000 1.8200
                 12.8800 1.8200 12.8800 0.9200 12.8850 0.9200 12.8850 0.8000 12.9750 0.8000
                 12.9750 0.5600 11.7050 0.5600 11.7050 1.1200 11.5650 1.1200 11.5650 0.8800
                 11.5850 0.8800 11.5850 0.4800 11.0650 0.4800 11.0650 1.1400 11.1850 1.1400
                 11.1850 1.2600 10.9450 1.2600 10.9450 0.9200 9.6450 0.9200 9.6450 1.1600 8.4050 1.1600
                 8.4050 1.0400 9.5250 1.0400 9.5250 0.8000 10.9450 0.8000 10.9450 0.3600 11.7050 0.3600
                 11.7050 0.4400 12.4050 0.4400 12.4050 0.3600 12.6450 0.3600 12.6450 0.4400
                 13.0950 0.4400 ;
        POLYGON  12.7650 0.8000 12.6450 0.8000 12.6450 1.4600 12.5650 1.4600 12.5650 1.8200
                 12.4450 1.8200 12.4450 1.4600 11.6650 1.4600 11.6650 2.2500 10.7600 2.2500
                 10.7600 1.7400 10.2800 1.7400 10.2800 2.0100 9.5600 2.0100 9.5600 1.6400 8.4450 1.6400
                 8.4450 2.0100 7.3650 2.0100 7.3650 1.0800 7.4850 1.0800 7.4850 1.8900 7.8450 1.8900
                 7.8450 0.9600 7.9250 0.9600 7.9250 0.8400 8.0450 0.8400 8.0450 1.0800 7.9650 1.0800
                 7.9650 1.8900 8.3250 1.8900 8.3250 1.5200 9.6800 1.5200 9.6800 1.8900 10.1600 1.8900
                 10.1600 1.6200 10.8800 1.6200 10.8800 2.1300 11.5450 2.1300 11.5450 1.2400
                 11.6650 1.2400 11.6650 1.3400 12.5250 1.3400 12.5250 0.6800 12.7650 0.6800 ;
        POLYGON  11.4650 0.7200 11.4250 0.7200 11.4250 1.6200 11.4050 1.6200 11.4050 2.0100
                 11.2850 2.0100 11.2850 1.5000 10.7050 1.5000 10.7050 1.1600 9.7650 1.1600
                 9.7650 1.0400 10.8250 1.0400 10.8250 1.3800 11.3050 1.3800 11.3050 0.7200
                 11.2250 0.7200 11.2250 0.6000 11.4650 0.6000 ;
        POLYGON  10.5850 1.4000 10.0400 1.4000 10.0400 1.7700 9.8000 1.7700 9.8000 1.6000 9.9200 1.6000
                 9.9200 1.4000 8.2050 1.4000 8.2050 1.7700 8.0850 1.7700 8.0850 1.2800 8.1650 1.2800
                 8.1650 0.5000 8.2850 0.5000 8.2850 0.7400 9.1650 0.7400 9.1650 0.6000 9.4050 0.6000
                 9.4050 0.7200 9.2850 0.7200 9.2850 0.8600 8.2850 0.8600 8.2850 1.2800 10.5850 1.2800 ;
        POLYGON  9.7650 0.6800 9.6450 0.6800 9.6450 0.4800 8.9850 0.4800 8.9850 0.6200 8.7450 0.6200
                 8.7450 0.5000 8.8650 0.5000 8.8650 0.3600 9.7650 0.3600 ;
        POLYGON  7.8650 0.7200 7.7250 0.7200 7.7250 1.7700 7.6050 1.7700 7.6050 0.9600 7.2450 0.9600
                 7.2450 1.1700 5.9850 1.1700 5.9850 0.9900 5.5050 0.9900 5.5050 0.5600 4.6850 0.5600
                 4.6850 0.5200 4.2750 0.5200 4.2750 1.2000 4.1550 1.2000 4.1550 0.4000 4.8050 0.4000
                 4.8050 0.4400 5.6250 0.4400 5.6250 0.8700 6.1050 0.8700 6.1050 1.0500 7.1250 1.0500
                 7.1250 0.8400 7.6050 0.8400 7.6050 0.6000 7.7450 0.6000 7.7450 0.4800 7.8650 0.4800 ;
        POLYGON  7.4850 0.6800 7.0050 0.6800 7.0050 0.9300 6.2250 0.9300 6.2250 0.7500 6.1050 0.7500
                 6.1050 0.6300 6.3450 0.6300 6.3450 0.8100 6.8850 0.8100 6.8850 0.5600 7.4850 0.5600 ;
        POLYGON  7.2450 1.6400 7.1250 1.6400 7.1250 1.5700 6.0650 1.5700 6.0650 1.7700 5.9450 1.7700
                 5.9450 1.4500 7.1250 1.4500 7.1250 1.4000 7.2450 1.4000 ;
        POLYGON  6.7650 0.6900 6.5250 0.6900 6.5250 0.5100 5.8650 0.5100 5.8650 0.7500 5.7450 0.7500
                 5.7450 0.3900 6.6450 0.3900 6.6450 0.5700 6.7650 0.5700 ;
        POLYGON  6.6050 2.2500 5.4650 2.2500 5.4650 1.6750 4.6850 1.6750 4.6850 0.6800 4.9650 0.6800
                 4.9650 0.8000 4.8050 0.8000 4.8050 1.5550 5.5850 1.5550 5.5850 2.1300 6.6050 2.1300 ;
        POLYGON  5.1050 2.2500 4.3350 2.2500 4.3350 1.8200 4.3950 1.8200 4.3950 1.4400 3.6150 1.4400
                 3.6150 2.2100 3.4950 2.2100 3.4950 1.2450 2.8750 1.2450 2.8750 1.1250 3.4950 1.1250
                 3.4950 0.6400 3.6150 0.6400 3.6150 1.3200 4.3950 1.3200 4.3950 0.6400 4.5150 0.6400
                 4.5150 1.9400 4.4550 1.9400 4.4550 2.1300 5.1050 2.1300 ;
    END
END DFFSRHQX8

MACRO DFFSRHQX4
    CLASS CORE ;
    FOREIGN DFFSRHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 0.5900 1.5150 1.9900 ;
        RECT  0.5550 1.0250 1.5150 1.1450 ;
        RECT  0.5550 0.8850 0.8000 1.1450 ;
        RECT  0.5550 0.5900 0.6750 1.9900 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9050 0.9400 3.1750 1.2000 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.1800 10.7150 1.4500 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6150 0.9400 11.8750 1.1550 ;
        RECT  11.6150 0.9400 11.7350 1.3200 ;
        END
    END CK
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2350 2.1300 8.4750 2.2500 ;
        RECT  7.5950 2.0100 8.3550 2.1300 ;
        RECT  7.5950 1.7000 7.7150 2.1300 ;
        RECT  6.9950 1.7000 7.7150 1.8200 ;
        RECT  5.7950 2.1300 7.1150 2.2500 ;
        RECT  6.9950 1.7000 7.1150 2.2500 ;
        RECT  5.7950 1.5200 5.9150 2.2500 ;
        RECT  5.2350 1.5200 5.9150 1.6400 ;
        RECT  5.2350 1.5200 5.4950 1.6700 ;
        RECT  5.0650 1.4300 5.3550 1.5500 ;
        END
    END SN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.8650 -0.1800 11.9850 0.8200 ;
        RECT  10.5150 -0.1800 10.6350 0.7800 ;
        RECT  9.1150 -0.1800 9.2350 0.6400 ;
        RECT  5.2050 -0.1800 5.4450 0.3400 ;
        RECT  2.5950 0.4600 2.8350 0.5800 ;
        RECT  2.7150 -0.1800 2.8350 0.5800 ;
        RECT  1.8150 -0.1800 1.9350 0.6400 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.8650 1.4600 11.9850 2.7900 ;
        RECT  10.6750 1.8400 10.7950 2.7900 ;
        RECT  8.5950 2.0100 8.8350 2.1300 ;
        RECT  8.5950 2.0100 8.7150 2.7900 ;
        RECT  7.3550 1.9400 7.4750 2.7900 ;
        RECT  7.2350 1.9400 7.4750 2.0600 ;
        RECT  5.0450 2.2700 5.2850 2.7900 ;
        RECT  3.7850 2.0400 3.9050 2.7900 ;
        RECT  3.6650 2.0400 3.9050 2.1600 ;
        RECT  2.6550 1.5600 2.7750 2.7900 ;
        RECT  1.8150 1.4400 1.9350 2.7900 ;
        RECT  0.9750 1.3400 1.0950 2.7900 ;
        RECT  0.1350 1.3400 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.6250 1.5600 11.3750 1.5600 11.3750 0.7000 11.4450 0.7000 11.4450 0.4800
                 10.8750 0.4800 10.8750 0.9400 11.0150 0.9400 11.0150 1.0600 10.7550 1.0600
                 10.7550 1.0400 10.1950 1.0400 10.1950 1.1600 10.0750 1.1600 10.0750 2.2500
                 9.4750 2.2500 9.4750 1.8900 7.8350 1.8900 7.8350 1.5800 6.8750 1.5800 6.8750 2.0100
                 6.2750 2.0100 6.2750 0.9800 6.3950 0.9800 6.3950 0.4900 5.9150 0.4900 5.9150 1.0700
                 5.6750 1.0700 5.6750 0.9500 5.7950 0.9500 5.7950 0.3700 6.5150 0.3700 6.5150 1.1000
                 6.3950 1.1000 6.3950 1.8900 6.7550 1.8900 6.7550 1.4600 7.9550 1.4600 7.9550 1.7700
                 9.4250 1.7700 9.4250 1.5400 9.3550 1.5400 9.3550 1.4200 9.5950 1.4200 9.5950 1.5400
                 9.5450 1.5400 9.5450 1.7700 9.5950 1.7700 9.5950 2.1300 9.9550 2.1300 9.9550 0.9200
                 10.7550 0.9200 10.7550 0.3600 11.5650 0.3600 11.5650 0.8200 11.4950 0.8200
                 11.4950 1.4400 11.6250 1.4400 ;
        POLYGON  11.2550 1.6900 11.2150 1.6900 11.2150 2.0800 11.0950 2.0800 11.0950 1.6900
                 10.1950 1.6900 10.1950 1.3400 10.3150 1.3400 10.3150 1.5700 11.1350 1.5700
                 11.1350 0.7200 10.9950 0.7200 10.9950 0.6000 11.2550 0.6000 ;
        POLYGON  9.9950 0.7400 9.8350 0.7400 9.8350 2.0100 9.7150 2.0100 9.7150 0.7400 9.4750 0.7400
                 9.4750 0.8800 8.7950 0.8800 8.7950 1.0000 8.5550 1.0000 8.5550 0.8800 8.6750 0.8800
                 8.6750 0.7600 9.3550 0.7600 9.3550 0.6200 9.8750 0.6200 9.8750 0.5000 9.9950 0.5000 ;
        POLYGON  9.5950 1.2400 8.3150 1.2400 8.3150 1.1000 6.8750 1.1000 6.8750 0.9800 8.4350 0.9800
                 8.4350 1.1200 9.3550 1.1200 9.3550 1.1000 9.5950 1.1000 ;
        POLYGON  9.2350 1.5400 8.3350 1.5400 8.3350 1.6500 8.0750 1.6500 8.0750 1.3400 6.6350 1.3400
                 6.6350 1.7700 6.5150 1.7700 6.5150 1.2200 6.6350 1.2200 6.6350 0.5500 6.7550 0.5500
                 6.7550 0.7400 7.8750 0.7400 7.8750 0.6000 8.1150 0.6000 8.1150 0.7200 7.9950 0.7200
                 7.9950 0.8600 6.7550 0.8600 6.7550 1.2200 8.1950 1.2200 8.1950 1.4200 9.2350 1.4200 ;
        POLYGON  8.4750 0.6800 8.3550 0.6800 8.3550 0.4800 7.7550 0.4800 7.7550 0.6200 7.4550 0.6200
                 7.4550 0.5000 7.6350 0.5000 7.6350 0.3600 8.4750 0.3600 ;
        POLYGON  6.2750 0.7300 6.1550 0.7300 6.1550 1.9700 6.0350 1.9700 6.0350 1.3100 4.9450 1.3100
                 4.9450 1.5700 4.4450 1.5700 4.4450 1.9200 2.8950 1.9200 2.8950 1.4400 2.5150 1.4400
                 2.5150 1.1200 2.6350 1.1200 2.6350 1.3200 3.0150 1.3200 3.0150 1.8000 4.3250 1.8000
                 4.3250 1.4500 4.8250 1.4500 4.8250 1.1900 6.0350 1.1900 6.0350 0.6100 6.2750 0.6100 ;
        POLYGON  5.6750 0.7300 5.4350 0.7300 5.4350 0.5800 4.9650 0.5800 4.9650 0.4800 4.4250 0.4800
                 4.4250 0.6200 4.1850 0.6200 4.1850 0.5000 4.3050 0.5000 4.3050 0.3600 5.0850 0.3600
                 5.0850 0.4600 5.5550 0.4600 5.5550 0.6100 5.6750 0.6100 ;
        POLYGON  5.6750 1.9100 4.6850 1.9100 4.6850 1.9700 4.5650 1.9700 4.5650 1.6900 4.6850 1.6900
                 4.6850 1.7900 5.6750 1.7900 ;
        POLYGON  5.6750 2.2500 5.4050 2.2500 5.4050 2.1500 4.9250 2.1500 4.9250 2.2100 4.7950 2.2100
                 4.7950 2.2500 4.0250 2.2500 4.0250 2.1300 4.6750 2.1300 4.6750 2.0900 4.8050 2.0900
                 4.8050 2.0300 5.5250 2.0300 5.5250 2.1300 5.6750 2.1300 ;
        POLYGON  4.8450 0.7200 4.7050 0.7200 4.7050 1.2800 3.7050 1.2800 3.7050 0.7200 3.5850 0.7200
                 3.5850 0.6000 3.8250 0.6000 3.8250 1.1600 4.5850 1.1600 4.5850 0.6000 4.8450 0.6000 ;
        POLYGON  4.4650 1.0400 4.2250 1.0400 4.2250 0.8600 3.9450 0.8600 3.9450 0.4800 3.0750 0.4800
                 3.0750 0.8200 2.3550 0.8200 2.3550 1.5600 2.4150 1.5600 2.4150 1.9000 2.1750 1.9000
                 2.1750 1.5600 2.2350 1.5600 2.2350 1.2000 1.6350 1.2000 1.6350 1.0800 2.2350 1.0800
                 2.2350 0.5000 2.3550 0.5000 2.3550 0.7000 2.9550 0.7000 2.9550 0.3600 4.0650 0.3600
                 4.0650 0.7400 4.3450 0.7400 4.3450 0.9200 4.4650 0.9200 ;
        POLYGON  3.5850 1.3000 3.4150 1.3000 3.4150 1.4400 3.2550 1.4400 3.2550 1.6800 3.1350 1.6800
                 3.1350 1.3200 3.2950 1.3200 3.2950 0.7200 3.1950 0.7200 3.1950 0.6000 3.4350 0.6000
                 3.4350 0.7200 3.4150 0.7200 3.4150 1.1800 3.5850 1.1800 ;
    END
END DFFSRHQX4

MACRO DFFSRHQX2
    CLASS CORE ;
    FOREIGN DFFSRHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0850 1.1000 2.3250 1.2900 ;
        RECT  2.1000 1.1000 2.2500 1.4700 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7250 2.1300 7.1850 2.2500 ;
        RECT  6.7250 1.7000 6.8450 2.2500 ;
        RECT  5.9250 1.7000 6.8450 1.8200 ;
        RECT  4.3050 2.1300 6.0450 2.2500 ;
        RECT  5.9250 1.7000 6.0450 2.2500 ;
        RECT  4.3050 1.6600 4.4250 2.2500 ;
        RECT  3.5200 1.6600 4.4250 1.7800 ;
        RECT  2.7250 1.8900 3.6400 2.0100 ;
        RECT  3.5200 1.6600 3.6400 2.0100 ;
        RECT  2.6250 1.2300 2.8850 1.3800 ;
        RECT  2.7250 1.1000 2.8450 2.0100 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2950 0.9400 9.5800 1.0900 ;
        RECT  9.1650 1.0800 9.4350 1.2000 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5100 0.8650 10.6600 1.3200 ;
        RECT  10.5100 0.8650 10.6300 1.3400 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.8100 0.8550 1.9600 ;
        RECT  0.5550 1.6000 0.7150 1.9600 ;
        RECT  0.5550 0.6800 0.6750 2.2100 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.7550 -0.1800 10.8750 0.7450 ;
        RECT  9.4050 -0.1800 9.6450 0.3400 ;
        RECT  7.8050 0.5000 8.0450 0.6200 ;
        RECT  7.8050 -0.1800 7.9250 0.6200 ;
        RECT  2.3450 0.6200 2.5850 0.7400 ;
        RECT  2.3450 -0.1800 2.4650 0.7400 ;
        RECT  0.9750 -0.1800 1.0950 0.8200 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.6900 1.4600 10.8100 2.7900 ;
        RECT  9.3850 1.5800 9.5050 2.7900 ;
        RECT  7.8050 2.0300 7.9250 2.7900 ;
        RECT  7.6850 2.0300 7.9250 2.1500 ;
        RECT  6.2850 1.9400 6.4050 2.7900 ;
        RECT  6.1650 1.9400 6.4050 2.0600 ;
        RECT  3.8250 1.9000 4.0650 2.0200 ;
        RECT  3.8250 1.9000 3.9450 2.7900 ;
        RECT  2.1250 1.8300 2.3650 1.9500 ;
        RECT  2.1650 1.8300 2.2850 2.7900 ;
        RECT  0.9750 1.6900 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.4550 0.7450 10.3900 0.7450 10.3900 1.5800 10.2700 1.5800 10.2700 0.5800
                 9.1750 0.5800 9.1750 0.9600 9.0450 0.9600 9.0450 1.1200 8.9250 1.1200 8.9250 0.8400
                 9.0550 0.8400 9.0550 0.4800 8.4250 0.4800 8.4250 1.2300 8.5450 1.2300 8.5450 1.3500
                 8.3050 1.3500 8.3050 0.8600 7.0050 0.8600 7.0050 1.1000 5.5650 1.1000 5.5650 0.9800
                 6.8850 0.9800 6.8850 0.7400 8.3050 0.7400 8.3050 0.3600 9.2850 0.3600 9.2850 0.4600
                 9.7650 0.4600 9.7650 0.3600 10.0050 0.3600 10.0050 0.4600 10.4550 0.4600 ;
        POLYGON  10.1250 0.8200 10.0050 0.8200 10.0050 1.4600 9.9250 1.4600 9.9250 1.8200 9.8050 1.8200
                 9.8050 1.4600 9.0250 1.4600 9.0250 2.2500 8.0450 2.2500 8.0450 1.9100 6.9650 1.9100
                 6.9650 1.5800 5.8050 1.5800 5.8050 2.0100 4.5450 2.0100 4.5450 1.2200 4.3850 1.2200
                 4.3850 1.1000 4.6650 1.1000 4.6650 1.8900 5.0250 1.8900 5.0250 0.8200 5.1450 0.8200
                 5.1450 1.8900 5.6850 1.8900 5.6850 1.4600 7.0850 1.4600 7.0850 1.7900 8.1650 1.7900
                 8.1650 2.1300 8.9050 2.1300 8.9050 1.2400 9.0250 1.2400 9.0250 1.3400 9.8850 1.3400
                 9.8850 0.7000 10.1250 0.7000 ;
        POLYGON  8.9350 0.7200 8.7850 0.7200 8.7850 1.7000 8.7650 1.7000 8.7650 2.0100 8.6450 2.0100
                 8.6450 1.5900 8.0650 1.5900 8.0650 1.1000 7.1250 1.1000 7.1250 0.9800 8.1850 0.9800
                 8.1850 1.4700 8.6650 1.4700 8.6650 0.6000 8.9350 0.6000 ;
        POLYGON  7.9450 1.3400 7.4450 1.3400 7.4450 1.6700 7.2050 1.6700 7.2050 1.5500 7.3250 1.5500
                 7.3250 1.3400 5.5650 1.3400 5.5650 1.7700 5.3250 1.7700 5.3250 0.7400 5.2650 0.7400
                 5.2650 0.5000 5.3850 0.5000 5.3850 0.6200 5.4450 0.6200 5.4450 0.7400 6.4650 0.7400
                 6.4650 0.6000 6.7650 0.6000 6.7650 0.7200 6.5850 0.7200 6.5850 0.8600 5.4450 0.8600
                 5.4450 1.2200 7.9450 1.2200 ;
        POLYGON  7.1850 0.6200 6.9450 0.6200 6.9450 0.4800 6.3450 0.4800 6.3450 0.6200 6.1050 0.6200
                 6.1050 0.5000 6.2250 0.5000 6.2250 0.3600 7.0650 0.3600 7.0650 0.5000 7.1850 0.5000 ;
        POLYGON  4.9050 1.7700 4.7850 1.7700 4.7850 0.9800 4.2650 0.9800 4.2650 1.2200 3.0050 1.2200
                 3.0050 0.9800 2.1050 0.9800 2.1050 0.4800 1.3350 0.4800 1.3350 1.2400 1.2150 1.2400
                 1.2150 0.3600 2.2250 0.3600 2.2250 0.8600 3.1250 0.8600 3.1250 1.1000 4.1450 1.1000
                 4.1450 0.8600 4.7850 0.8600 4.7850 0.5000 4.9050 0.5000 ;
        POLYGON  4.5450 0.6800 4.4250 0.6800 4.4250 0.7400 4.0250 0.7400 4.0250 0.9800 3.3050 0.9800
                 3.3050 0.7400 3.1850 0.7400 3.1850 0.6200 3.4250 0.6200 3.4250 0.8600 3.9050 0.8600
                 3.9050 0.6200 4.3050 0.6200 4.3050 0.5600 4.5450 0.5600 ;
        POLYGON  4.4250 1.5400 3.2050 1.5400 3.2050 1.7700 2.9650 1.7700 2.9650 1.5300 3.0850 1.5300
                 3.0850 1.4200 4.4250 1.4200 ;
        POLYGON  3.7850 0.7400 3.6650 0.7400 3.6650 0.5000 2.9450 0.5000 2.9450 0.7400 2.8250 0.7400
                 2.8250 0.3800 3.7850 0.3800 ;
        POLYGON  3.7050 2.2500 2.4850 2.2500 2.4850 1.7100 1.7050 1.7100 1.7050 0.7200 1.8650 0.7200
                 1.8650 0.6000 1.9850 0.6000 1.9850 0.8400 1.8250 0.8400 1.8250 1.5900 2.6050 1.5900
                 2.6050 2.1300 3.7050 2.1300 ;
        POLYGON  2.0450 2.2500 1.3950 2.2500 1.3950 1.8000 1.4550 1.8000 1.4550 1.4800 0.8150 1.4800
                 0.8150 1.2200 0.9350 1.2200 0.9350 1.3600 1.4550 1.3600 1.4550 0.6800 1.5750 0.6800
                 1.5750 1.9200 1.5150 1.9200 1.5150 2.1300 2.0450 2.1300 ;
    END
END DFFSRHQX2

MACRO DFFSRHQX1
    CLASS CORE ;
    FOREIGN DFFSRHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7250 1.1900 2.0150 1.3800 ;
        RECT  1.6550 1.1700 1.9250 1.3300 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9700 2.1300 6.4750 2.2500 ;
        RECT  5.9700 1.7600 6.0900 2.2500 ;
        RECT  5.2150 1.7600 6.0900 1.8800 ;
        RECT  3.7450 2.1300 5.3350 2.2500 ;
        RECT  5.2150 1.7600 5.3350 2.2500 ;
        RECT  3.7450 1.7000 3.8650 2.2500 ;
        RECT  3.1000 1.7000 3.8650 1.8200 ;
        RECT  2.3050 1.8900 3.2200 2.0100 ;
        RECT  3.1000 1.7000 3.2200 2.0100 ;
        RECT  2.3050 1.1750 2.5400 1.4350 ;
        RECT  2.2550 1.1700 2.4950 1.2900 ;
        RECT  2.3050 1.1700 2.4250 2.0100 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5750 1.2300 8.9750 1.3800 ;
        RECT  8.5750 1.2100 8.7150 1.4500 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.8750 1.1750 10.1350 1.3800 ;
        RECT  9.8750 1.0300 9.9950 1.3800 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  10.1150 -0.1800 10.2350 0.9100 ;
        RECT  8.7350 -0.1800 8.8550 0.8500 ;
        RECT  7.1550 -0.1800 7.2750 0.6800 ;
        RECT  1.9750 -0.1800 2.0950 0.8100 ;
        RECT  0.5550 -0.1800 0.6750 0.8200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  10.1150 1.5000 10.2350 2.7900 ;
        RECT  8.6750 1.8100 8.7950 2.7900 ;
        RECT  7.2150 1.9300 7.3350 2.7900 ;
        RECT  7.0950 1.9300 7.3350 2.0500 ;
        RECT  5.5750 2.0000 5.6950 2.7900 ;
        RECT  5.4550 2.0000 5.6950 2.1200 ;
        RECT  3.3850 1.9400 3.6250 2.0600 ;
        RECT  3.3850 1.9400 3.5050 2.7900 ;
        RECT  1.8250 1.7400 1.9450 2.7900 ;
        RECT  1.7050 1.7400 1.9450 1.8600 ;
        RECT  0.5550 1.6900 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.8750 1.6200 9.6350 1.6200 9.6350 0.7900 9.6950 0.7900 9.6950 0.5600 9.0950 0.5600
                 9.0950 1.0900 8.4550 1.0900 8.4550 1.1300 8.1950 1.1300 8.1950 1.0100 8.3350 1.0100
                 8.3350 0.4800 7.7150 0.4800 7.7150 1.2100 7.8350 1.2100 7.8350 1.3300 7.5950 1.3300
                 7.5950 0.9200 6.2950 0.9200 6.2950 1.1600 5.0350 1.1600 5.0350 1.0400 6.1750 1.0400
                 6.1750 0.8000 7.5950 0.8000 7.5950 0.3600 8.4550 0.3600 8.4550 0.9700 8.9750 0.9700
                 8.9750 0.4400 9.0150 0.4400 9.0150 0.3600 9.2550 0.3600 9.2550 0.4400 9.8150 0.4400
                 9.8150 0.9100 9.7550 0.9100 9.7550 1.5000 9.8750 1.5000 ;
        POLYGON  9.4550 1.3300 9.2150 1.3300 9.2150 2.0500 9.0950 2.0500 9.0950 1.6900 8.3150 1.6900
                 8.3150 2.2500 7.4550 2.2500 7.4550 1.8100 6.9750 1.8100 6.9750 2.0100 6.2550 2.0100
                 6.2550 1.6400 5.0950 1.6400 5.0950 2.0100 4.0150 2.0100 4.0150 1.0600 4.1350 1.0600
                 4.1350 1.8900 4.4950 1.8900 4.4950 1.0400 4.5550 1.0400 4.5550 0.8400 4.6750 0.8400
                 4.6750 1.1600 4.6150 1.1600 4.6150 1.8900 4.9750 1.8900 4.9750 1.5200 6.3750 1.5200
                 6.3750 1.8900 6.8550 1.8900 6.8550 1.6900 7.5750 1.6900 7.5750 2.1300 8.1950 2.1300
                 8.1950 1.3100 8.3150 1.3100 8.3150 1.5700 9.0950 1.5700 9.0950 1.2100 9.2150 1.2100
                 9.2150 0.6800 9.4550 0.6800 ;
        POLYGON  8.2150 0.7200 8.0750 0.7200 8.0750 1.6900 8.0550 1.6900 8.0550 2.0100 7.9350 2.0100
                 7.9350 1.5700 7.3550 1.5700 7.3550 1.1600 6.4150 1.1600 6.4150 1.0400 7.4750 1.0400
                 7.4750 1.4500 7.9550 1.4500 7.9550 0.6000 8.2150 0.6000 ;
        POLYGON  7.2350 1.4000 6.7350 1.4000 6.7350 1.7700 6.4950 1.7700 6.4950 1.6500 6.6150 1.6500
                 6.6150 1.4000 4.8550 1.4000 4.8550 1.7700 4.7350 1.7700 4.7350 1.2800 4.7950 1.2800
                 4.7950 0.5000 4.9150 0.5000 4.9150 0.7400 5.8150 0.7400 5.8150 0.6000 6.0550 0.6000
                 6.0550 0.7200 5.9350 0.7200 5.9350 0.8600 4.9150 0.8600 4.9150 1.2800 7.2350 1.2800 ;
        POLYGON  6.4150 0.6800 6.2950 0.6800 6.2950 0.4800 5.6350 0.4800 5.6350 0.6200 5.3950 0.6200
                 5.3950 0.5000 5.5150 0.5000 5.5150 0.3600 6.4150 0.3600 ;
        POLYGON  4.4350 0.9200 4.3750 0.9200 4.3750 1.7700 4.2550 1.7700 4.2550 0.9400 3.8950 0.9400
                 3.8950 1.2300 2.6600 1.2300 2.6600 1.0500 1.7350 1.0500 1.7350 0.5100 0.9150 0.5100
                 0.9150 1.2400 0.7950 1.2400 0.7950 0.3900 1.8550 0.3900 1.8550 0.9300 2.7800 0.9300
                 2.7800 1.1100 3.7750 1.1100 3.7750 0.8200 4.2550 0.8200 4.2550 0.8000 4.3150 0.8000
                 4.3150 0.5000 4.4350 0.5000 ;
        POLYGON  4.0750 0.6800 3.9550 0.6800 3.9550 0.7000 3.6550 0.7000 3.6550 0.9900 2.9000 0.9900
                 2.9000 0.8100 2.7550 0.8100 2.7550 0.6900 3.0200 0.6900 3.0200 0.8700 3.5350 0.8700
                 3.5350 0.5800 3.8350 0.5800 3.8350 0.5600 4.0750 0.5600 ;
        POLYGON  3.8950 1.5800 2.7850 1.5800 2.7850 1.7700 2.5450 1.7700 2.5450 1.5550 2.6650 1.5550
                 2.6650 1.4600 3.8950 1.4600 ;
        POLYGON  3.4150 0.7500 3.1750 0.7500 3.1750 0.5700 2.5150 0.5700 2.5150 0.8100 2.3950 0.8100
                 2.3950 0.4500 3.2950 0.4500 3.2950 0.6300 3.4150 0.6300 ;
        POLYGON  3.2650 2.2500 2.0650 2.2500 2.0650 1.6200 1.4050 1.6200 1.4050 1.6700 1.2850 1.6700
                 1.2850 0.6300 1.6150 0.6300 1.6150 0.7500 1.4050 0.7500 1.4050 1.5000 2.1850 1.5000
                 2.1850 2.1300 3.2650 2.1300 ;
        POLYGON  1.7050 2.2500 0.9750 2.2500 0.9750 1.8200 1.0350 1.8200 1.0350 1.4800 0.4150 1.4800
                 0.4150 1.2400 0.5350 1.2400 0.5350 1.3600 1.0350 1.3600 1.0350 0.6800 1.1550 0.6800
                 1.1550 1.9400 1.0950 1.9400 1.0950 2.1300 1.7050 2.1300 ;
    END
END DFFSRHQX1

MACRO DFFSHQX8
    CLASS CORE ;
    FOREIGN DFFSHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7900 0.6550 2.9100 2.2100 ;
        RECT  0.0700 1.0250 2.9100 1.1450 ;
        RECT  1.9500 0.6550 2.0700 2.2100 ;
        RECT  1.1100 0.6550 1.2300 2.2050 ;
        RECT  0.2700 0.6550 0.3900 2.2050 ;
        RECT  0.0700 0.8850 0.3900 1.1450 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8400 0.4900 7.9600 1.2300 ;
        RECT  7.3400 0.4900 7.9600 0.6100 ;
        RECT  7.3400 0.3600 7.4600 0.6100 ;
        RECT  5.5800 0.3600 7.4600 0.4800 ;
        RECT  5.5800 0.8850 5.7300 1.1450 ;
        RECT  5.5800 0.3600 5.7000 1.3400 ;
        RECT  5.1600 1.2200 5.7000 1.3400 ;
        RECT  5.0400 1.2600 5.2800 1.3800 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.1600 1.1400 10.4250 1.3850 ;
        RECT  10.1650 1.1200 10.4250 1.3850 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.6000 1.2100 11.0050 1.3850 ;
        RECT  10.7450 1.1800 11.0050 1.3850 ;
        END
    END CK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.4000 -0.1800 10.5200 0.7400 ;
        RECT  8.8200 0.4600 9.0600 0.5800 ;
        RECT  8.8200 -0.1800 8.9400 0.5800 ;
        RECT  7.5800 -0.1800 7.8200 0.3700 ;
        RECT  4.8400 -0.1800 4.9600 0.6800 ;
        RECT  4.0000 -0.1800 4.1200 0.7300 ;
        RECT  3.2700 -0.1800 3.3900 0.5300 ;
        RECT  2.3700 -0.1800 2.4900 0.6450 ;
        RECT  1.5300 -0.1800 1.6500 0.6450 ;
        RECT  0.6900 -0.1800 0.8100 0.6450 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.2800 1.7450 10.4000 2.7900 ;
        RECT  8.8800 2.0700 9.0000 2.7900 ;
        RECT  8.7600 2.0700 9.0000 2.1900 ;
        RECT  8.1600 2.2900 8.4000 2.7900 ;
        RECT  5.6200 1.9800 5.8600 2.1500 ;
        RECT  5.6200 1.9800 5.7400 2.7900 ;
        RECT  4.8400 1.7400 4.9600 2.7900 ;
        RECT  4.0000 1.5600 4.1200 2.7900 ;
        RECT  3.2100 1.9700 3.3300 2.7900 ;
        RECT  2.3700 1.4650 2.4900 2.7900 ;
        RECT  1.5300 1.4650 1.6500 2.7900 ;
        RECT  0.6900 1.4650 0.8100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.9400 0.7400 10.7600 0.7400 10.7600 1.0000 10.0400 1.0000 10.0400 1.5050
                 10.8200 1.5050 10.8200 1.9000 10.7000 1.9000 10.7000 1.6250 10.0400 1.6250
                 10.0400 2.2300 9.5600 2.2300 9.5600 2.2500 9.3200 2.2500 9.3200 2.1300 9.3600 2.1300
                 9.3600 1.9500 8.6400 1.9500 8.6400 2.0700 8.3750 2.0700 8.3750 2.1700 8.0400 2.1700
                 8.0400 2.2500 7.4800 2.2500 7.4800 2.1300 7.9200 2.1300 7.9200 2.0500 8.2550 2.0500
                 8.2550 1.9500 8.5200 1.9500 8.5200 1.8300 9.4800 1.8300 9.4800 2.1100 9.9200 2.1100
                 9.9200 1.0000 9.8400 1.0000 9.8400 0.8800 10.6400 0.8800 10.6400 0.6200 10.8200 0.6200
                 10.8200 0.5000 10.9400 0.5000 ;
        POLYGON  9.7400 0.7600 9.7200 0.7600 9.7200 1.9900 9.6000 1.9900 9.6000 1.3300 8.5600 1.3300
                 8.5600 1.2100 9.6000 1.2100 9.6000 0.6400 9.6200 0.6400 9.6200 0.5000 9.7400 0.5000 ;
        POLYGON  9.4800 1.0800 9.3600 1.0800 9.3600 0.8400 8.5800 0.8400 8.5800 0.5500 8.2000 0.5500
                 8.2000 1.4700 7.4400 1.4700 7.4400 1.6500 7.5600 1.6500 7.5600 1.7700 7.3200 1.7700
                 7.3200 0.9000 6.6200 0.9000 6.6200 0.6600 6.7400 0.6600 6.7400 0.7800 7.1000 0.7800
                 7.1000 0.7300 7.3400 0.7300 7.3400 0.7800 7.4400 0.7800 7.4400 1.3500 8.0800 1.3500
                 8.0800 0.4300 8.7000 0.4300 8.7000 0.7200 9.4800 0.7200 ;
        POLYGON  9.2200 1.0900 8.4400 1.0900 8.4400 1.4700 8.4600 1.4700 8.4600 1.7100 8.4000 1.7100
                 8.4000 1.8300 7.8000 1.8300 7.8000 2.0100 7.1100 2.0100 7.1100 2.2100 6.9900 2.2100
                 6.9900 1.6900 7.0100 1.6900 7.0100 1.1400 6.3800 1.1400 6.3800 0.7200 6.2400 0.7200
                 6.2400 0.6000 6.5000 0.6000 6.5000 1.0200 7.1300 1.0200 7.1300 1.8900 7.6800 1.8900
                 7.6800 1.7100 8.2800 1.7100 8.2800 1.5900 8.3200 1.5900 8.3200 0.7900 8.3400 0.7900
                 8.3400 0.6700 8.4600 0.6700 8.4600 0.9700 9.2200 0.9700 ;
        POLYGON  6.8900 1.3800 6.0900 1.3800 6.0900 1.1000 6.2100 1.1000 6.2100 1.2600 6.8900 1.2600 ;
        POLYGON  6.6900 2.2100 6.5700 2.2100 6.5700 1.6200 4.8000 1.6200 4.8000 1.4200 4.6400 1.4200
                 4.6400 1.3000 4.9200 1.3000 4.9200 1.5000 5.8500 1.5000 5.8500 0.7200 5.8200 0.7200
                 5.8200 0.6000 6.0600 0.6000 6.0600 0.7200 5.9700 0.7200 5.9700 1.5000 6.6900 1.5000 ;
        POLYGON  6.2700 2.2100 6.1500 2.2100 6.1500 1.8600 5.3800 1.8600 5.3800 2.2100 5.2600 2.2100
                 5.2600 1.7400 6.2700 1.7400 ;
        POLYGON  5.4600 1.1000 4.5200 1.1000 4.5200 1.5600 4.5400 1.5600 4.5400 2.2100 4.4200 2.2100
                 4.4200 1.6800 4.4000 1.6800 4.4000 1.1000 3.7000 1.1000 3.7000 1.8200 3.5800 1.8200
                 3.5800 1.1000 3.1900 1.1000 3.1900 1.2200 3.0700 1.2200 3.0700 0.9800 3.5800 0.9800
                 3.5800 0.6800 3.7000 0.6800 3.7000 0.9800 4.4000 0.9800 4.4000 0.8600 4.4200 0.8600
                 4.4200 0.6300 4.5400 0.6300 4.5400 0.9800 5.3400 0.9800 5.3400 0.8600 5.4600 0.8600 ;
    END
END DFFSHQX8

MACRO DFFSHQX4
    CLASS CORE ;
    FOREIGN DFFSHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 0.6300 1.6700 2.2100 ;
        RECT  0.6500 1.3150 1.6700 1.4350 ;
        RECT  0.7100 0.6300 0.8300 2.2100 ;
        RECT  0.6500 1.1750 0.8300 1.4350 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.4850 0.7000 5.6050 1.0800 ;
        RECT  4.9550 0.7000 5.6050 0.8200 ;
        RECT  4.9550 0.3600 5.0750 0.8200 ;
        RECT  3.8950 0.3600 5.0750 0.4800 ;
        RECT  3.5500 0.4400 4.0150 0.5600 ;
        RECT  3.5500 0.8850 3.7000 1.1450 ;
        RECT  2.9100 1.2200 3.6700 1.3400 ;
        RECT  3.5500 0.4400 3.6700 1.3400 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8450 1.1800 8.1050 1.4100 ;
        RECT  7.9050 1.0200 8.0250 1.4300 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.2150 1.0200 9.3350 1.2600 ;
        RECT  9.0050 1.2300 9.2650 1.3800 ;
        RECT  9.1450 1.1400 9.3350 1.2600 ;
        END
    END CK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.4550 -0.1800 9.5750 0.9200 ;
        RECT  7.9250 0.5400 8.1650 0.6600 ;
        RECT  7.9250 -0.1800 8.0450 0.6600 ;
        RECT  6.4050 -0.1800 6.5250 0.6900 ;
        RECT  5.2650 0.4600 5.5050 0.5800 ;
        RECT  5.3850 -0.1800 5.5050 0.5800 ;
        RECT  2.8100 -0.1800 2.9300 0.6800 ;
        RECT  1.9700 -0.1800 2.0900 0.6800 ;
        RECT  1.1300 -0.1800 1.2500 0.6800 ;
        RECT  0.2900 -0.1800 0.4100 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  9.3950 1.4600 9.5150 2.7900 ;
        RECT  8.0650 1.7900 8.1850 2.7900 ;
        RECT  6.3100 2.2900 6.5500 2.7900 ;
        RECT  5.3500 2.2900 5.5900 2.7900 ;
        RECT  3.6500 1.9400 3.7700 2.7900 ;
        RECT  2.8100 1.7000 2.9300 2.7900 ;
        RECT  1.9700 1.6900 2.0900 2.7900 ;
        RECT  1.1300 1.5600 1.2500 2.7900 ;
        RECT  0.2900 1.5600 0.4100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.1550 1.6200 8.7650 1.6200 8.7650 0.8400 8.9750 0.8400 8.9750 0.4800 8.4050 0.4800
                 8.4050 1.0600 8.1650 1.0600 8.1650 0.9000 7.6650 0.9000 7.6650 1.0500 7.4450 1.0500
                 7.4450 1.9300 5.2050 1.9300 5.2050 1.8600 4.8600 1.8600 4.8600 1.3000 4.1800 1.3000
                 4.1800 1.0400 4.0600 1.0400 4.0600 0.9200 4.3000 0.9200 4.3000 1.1800 5.1000 1.1800
                 5.1000 1.3000 4.9800 1.3000 4.9800 1.7400 5.3250 1.7400 5.3250 1.8100 7.3250 1.8100
                 7.3250 1.2900 6.8450 1.2900 6.8450 1.1700 7.3250 1.1700 7.3250 0.7800 8.2850 0.7800
                 8.2850 0.3600 9.0950 0.3600 9.0950 0.9600 8.8850 0.9600 8.8850 1.5000 9.1550 1.5000 ;
        POLYGON  8.7650 0.7200 8.6450 0.7200 8.6450 1.3000 8.6050 1.3000 8.6050 1.9100 8.4850 1.9100
                 8.4850 1.6700 7.6850 1.6700 7.6850 2.1700 5.1700 2.1700 5.1700 2.2400 4.4000 2.2400
                 4.4000 2.1200 5.0500 2.1200 5.0500 2.0500 7.5650 2.0500 7.5650 1.1900 7.6850 1.1900
                 7.6850 1.5500 8.4850 1.5500 8.4850 1.1800 8.5250 1.1800 8.5250 0.6000 8.7650 0.6000 ;
        POLYGON  7.5250 0.6600 7.2050 0.6600 7.2050 1.0500 6.7250 1.0500 6.7250 1.4500 7.0850 1.4500
                 7.0850 1.5700 7.2050 1.5700 7.2050 1.6900 6.9650 1.6900 6.9650 1.5700 6.6050 1.5700
                 6.6050 1.2900 6.0850 1.2900 6.0850 1.3300 5.9650 1.3300 5.9650 1.0900 6.0850 1.0900
                 6.0850 1.1700 6.6050 1.1700 6.6050 0.9300 7.0850 0.9300 7.0850 0.5400 7.5250 0.5400 ;
        POLYGON  6.4850 1.0500 6.2050 1.0500 6.2050 0.9700 5.8450 0.9700 5.8450 1.5700 6.0700 1.5700
                 6.0700 1.6900 5.7250 1.6900 5.7250 1.3200 5.3400 1.3200 5.3400 1.6200 5.1000 1.6200
                 5.1000 1.5000 5.2200 1.5000 5.2200 1.0600 4.7150 1.0600 4.7150 0.7200 4.5600 0.7200
                 4.5600 0.6000 4.8350 0.6000 4.8350 0.9400 5.3400 0.9400 5.3400 1.2000 5.7250 1.2000
                 5.7250 0.8500 5.9650 0.8500 5.9650 0.5000 6.0850 0.5000 6.0850 0.8500 6.3250 0.8500
                 6.3250 0.9300 6.4850 0.9300 ;
        POLYGON  4.7400 1.9600 4.6200 1.9600 4.6200 1.5800 2.6300 1.5800 2.6300 1.3300 2.7500 1.3300
                 2.7500 1.4600 3.8200 1.4600 3.8200 0.6800 4.1400 0.6800 4.1400 0.6000 4.3800 0.6000
                 4.3800 0.7200 4.2600 0.7200 4.2600 0.8000 3.9400 0.8000 3.9400 1.4600 4.6200 1.4600
                 4.6200 1.4400 4.7400 1.4400 ;
        POLYGON  4.3800 1.9000 4.1400 1.9000 4.1400 1.8200 3.3500 1.8200 3.3500 2.2100 3.2300 2.2100
                 3.2300 1.7000 4.3800 1.7000 ;
        POLYGON  3.4300 1.1000 3.3100 1.1000 3.3100 1.0700 2.5100 1.0700 2.5100 2.2100 2.3900 2.2100
                 2.3900 1.0700 1.9500 1.0700 1.9500 1.1900 1.8300 1.1900 1.8300 0.9500 2.3900 0.9500
                 2.3900 0.5400 2.5100 0.5400 2.5100 0.9500 3.3100 0.9500 3.3100 0.8600 3.4300 0.8600 ;
    END
END DFFSHQX4

MACRO DFFSHQX2
    CLASS CORE ;
    FOREIGN DFFSHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9800 0.8800 5.1000 1.2400 ;
        RECT  4.6100 0.8800 5.1000 1.0000 ;
        RECT  4.6100 0.3600 4.7300 1.0000 ;
        RECT  2.6800 0.3600 4.7300 0.4800 ;
        RECT  2.6800 0.8850 2.8300 1.1450 ;
        RECT  2.6800 0.3600 2.8000 1.3400 ;
        RECT  2.2600 1.2200 2.8000 1.3400 ;
        RECT  2.1400 1.2600 2.3800 1.3800 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 1.1200 7.5250 1.3900 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8450 1.1650 8.1050 1.3900 ;
        RECT  7.7200 1.1650 8.1050 1.3650 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 0.6400 0.8000 1.9900 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.5200 -0.1800 7.6400 0.7400 ;
        RECT  5.8800 -0.1800 6.1200 0.3200 ;
        RECT  4.8500 0.6400 5.0900 0.7600 ;
        RECT  4.8500 -0.1800 4.9700 0.7600 ;
        RECT  1.9400 -0.1800 2.0600 0.6800 ;
        RECT  1.1000 -0.1800 1.2200 0.6900 ;
        RECT  0.2600 -0.1800 0.3800 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.4000 1.7500 7.5200 2.7900 ;
        RECT  6.0600 1.6800 6.1800 2.7900 ;
        RECT  5.9400 1.6800 6.1800 1.9300 ;
        RECT  4.9200 2.2900 5.1600 2.7900 ;
        RECT  2.7200 1.9800 2.9600 2.1500 ;
        RECT  2.7200 1.9800 2.8400 2.7900 ;
        RECT  1.9400 1.7400 2.0600 2.7900 ;
        RECT  1.1000 1.3400 1.2200 2.7900 ;
        RECT  0.2600 1.3400 0.3800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.0600 1.0000 7.1450 1.0000 7.1450 1.5100 7.8100 1.5100 7.8100 1.6600 7.9400 1.6600
                 7.9400 1.9000 7.8200 1.9000 7.8200 1.7800 7.6900 1.7800 7.6900 1.6300 7.2800 1.6300
                 7.2800 2.2300 6.6800 2.2300 6.6800 2.2500 6.4400 2.2500 6.4400 2.1300 6.4800 2.1300
                 6.4800 1.5600 5.8200 1.5600 5.8200 2.1700 4.6000 2.1700 4.6000 2.0500 5.7000 2.0500
                 5.7000 1.4400 6.6000 1.4400 6.6000 2.1100 7.0250 2.1100 7.0250 1.0000 6.9600 1.0000
                 6.9600 0.8800 7.9400 0.8800 7.9400 0.5000 8.0600 0.5000 ;
        POLYGON  6.8600 0.7600 6.8400 0.7600 6.8400 1.9900 6.7200 1.9900 6.7200 1.3200 5.7000 1.3200
                 5.7000 1.2000 6.7200 1.2000 6.7200 0.6400 6.7400 0.6400 6.7400 0.5000 6.8600 0.5000 ;
        POLYGON  6.6000 1.0800 6.4800 1.0800 6.4800 0.8400 6.2150 0.8400 6.2150 0.5600 5.3400 0.5600
                 5.3400 1.4800 4.6600 1.4800 4.6600 1.6900 4.3700 1.6900 4.3700 1.1400 4.2300 1.1400
                 4.2300 0.9000 4.3700 0.9000 4.3700 0.7600 4.2500 0.7600 4.2500 0.6400 4.4900 0.6400
                 4.4900 1.3600 5.2200 1.3600 5.2200 0.4400 6.3350 0.4400 6.3350 0.7200 6.6000 0.7200 ;
        POLYGON  6.3400 1.0800 5.5800 1.0800 5.5800 1.9300 4.2100 1.9300 4.2100 2.2100 4.0900 2.2100
                 4.0900 1.3800 3.9900 1.3800 3.9900 0.7200 3.6100 0.7200 3.6100 0.6000 4.1100 0.6000
                 4.1100 1.2600 4.2100 1.2600 4.2100 1.8100 5.4600 1.8100 5.4600 0.9600 5.5500 0.9600
                 5.5500 0.6800 5.6700 0.6800 5.6700 0.9600 6.3400 0.9600 ;
        POLYGON  3.8700 1.3600 3.7500 1.3600 3.7500 1.2400 3.1900 1.2400 3.1900 0.8800 3.3100 0.8800
                 3.3100 1.1200 3.8700 1.1200 ;
        POLYGON  3.7900 2.2100 3.6700 2.2100 3.6700 1.6000 3.0700 1.6000 3.0700 1.6200 1.8000 1.6200
                 1.8000 1.3700 1.9200 1.3700 1.9200 1.5000 2.9500 1.5000 2.9500 0.6400 3.1900 0.6400
                 3.1900 0.6000 3.4300 0.6000 3.4300 0.7200 3.3100 0.7200 3.3100 0.7600 3.0700 0.7600
                 3.0700 1.4800 3.7900 1.4800 ;
        POLYGON  3.3700 2.2100 3.2500 2.2100 3.2500 1.8600 2.4800 1.8600 2.4800 2.2100 2.3600 2.2100
                 2.3600 1.7400 3.2500 1.7400 3.2500 1.7200 3.3700 1.7200 ;
        POLYGON  2.5600 1.1000 1.6400 1.1000 1.6400 2.2100 1.5200 2.2100 1.5200 1.1000 1.0600 1.1000
                 1.0600 1.2200 0.9400 1.2200 0.9400 0.9800 1.5200 0.9800 1.5200 0.5400 1.6400 0.5400
                 1.6400 0.9800 2.4400 0.9800 2.4400 0.8600 2.5600 0.8600 ;
    END
END DFFSHQX2

MACRO DFFSHQX1
    CLASS CORE ;
    FOREIGN DFFSHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6350 0.8500 4.7550 1.1500 ;
        RECT  4.2350 0.8500 4.7550 0.9700 ;
        RECT  4.2350 0.3600 4.3550 0.9700 ;
        RECT  2.3900 0.3600 4.3550 0.4800 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.3900 0.3600 2.5100 1.3400 ;
        RECT  1.9700 1.2200 2.5100 1.3400 ;
        RECT  1.8500 1.2600 2.0900 1.3800 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9750 1.1200 7.2350 1.3900 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5550 1.1650 7.8150 1.3800 ;
        RECT  7.4350 1.1200 7.6750 1.3100 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4200 0.6400 0.5400 1.9900 ;
        RECT  0.0700 1.1750 0.5400 1.2950 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.2950 -0.1800 7.4150 0.7400 ;
        RECT  5.7150 0.4600 5.9550 0.5800 ;
        RECT  5.7150 -0.1800 5.8350 0.5800 ;
        RECT  4.4750 0.6100 4.7150 0.7300 ;
        RECT  4.4750 -0.1800 4.5950 0.7300 ;
        RECT  1.6500 -0.1800 1.7700 0.6800 ;
        RECT  0.8400 -0.1800 0.9600 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.0950 1.7500 7.2150 2.7900 ;
        RECT  5.7350 1.6800 5.8550 2.7900 ;
        RECT  4.6550 2.2300 4.8950 2.7900 ;
        RECT  2.4300 1.9800 2.6700 2.1500 ;
        RECT  2.4300 1.9800 2.5500 2.7900 ;
        RECT  1.6500 1.7400 1.7700 2.7900 ;
        RECT  0.8400 1.3400 0.9600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.8350 0.8800 7.6550 0.8800 7.6550 1.0000 6.8550 1.0000 6.8550 1.5100 7.5050 1.5100
                 7.5050 1.6600 7.6350 1.6600 7.6350 1.9000 7.5150 1.9000 7.5150 1.7800 7.3850 1.7800
                 7.3850 1.6300 6.9750 1.6300 6.9750 2.2100 6.3950 2.2100 6.3950 2.2500 6.1550 2.2500
                 6.1550 2.1300 6.2050 2.1300 6.2050 1.5600 5.6150 1.5600 5.6150 2.2100 5.0150 2.2100
                 5.0150 2.1100 4.3350 2.1100 4.3350 1.9900 5.1350 1.9900 5.1350 2.0900 5.4950 2.0900
                 5.4950 1.4400 6.3250 1.4400 6.3250 2.0900 6.7350 2.0900 6.7350 0.8800 7.5350 0.8800
                 7.5350 0.7600 7.7150 0.7600 7.7150 0.5000 7.8350 0.5000 ;
        POLYGON  6.6350 0.7600 6.6150 0.7600 6.6150 1.3200 6.5750 1.3200 6.5750 1.9700 6.4550 1.9700
                 6.4550 1.3200 5.4750 1.3200 5.4750 1.1900 5.7150 1.1900 5.7150 1.2000 6.4950 1.2000
                 6.4950 0.6400 6.5150 0.6400 6.5150 0.5000 6.6350 0.5000 ;
        POLYGON  6.3750 1.0800 6.2550 1.0800 6.2550 0.8300 5.4750 0.8300 5.4750 0.5300 4.9950 0.5300
                 4.9950 1.3900 4.2950 1.3900 4.2950 1.5100 4.4150 1.5100 4.4150 1.6300 4.1750 1.6300
                 4.1750 1.2100 3.9800 1.2100 3.9800 0.7300 3.8750 0.7300 3.8750 0.6100 4.1150 0.6100
                 4.1150 0.7300 4.1000 0.7300 4.1000 1.0900 4.2950 1.0900 4.2950 1.2700 4.8750 1.2700
                 4.8750 0.4100 5.5950 0.4100 5.5950 0.7100 6.3750 0.7100 ;
        POLYGON  6.0750 1.0700 5.3550 1.0700 5.3550 1.4500 5.3750 1.4500 5.3750 1.9700 5.2550 1.9700
                 5.2550 1.8700 3.9200 1.8700 3.9200 2.2100 3.8000 2.2100 3.8000 1.4500 3.7400 1.4500
                 3.7400 0.9700 3.0500 0.9700 3.0500 0.6000 3.2900 0.6000 3.2900 0.8500 3.8600 0.8500
                 3.8600 1.3300 3.9200 1.3300 3.9200 1.7500 5.2550 1.7500 5.2550 1.5700 5.2350 1.5700
                 5.2350 0.7700 5.1150 0.7700 5.1150 0.6500 5.3550 0.6500 5.3550 0.9500 6.0750 0.9500 ;
        POLYGON  3.6200 1.3400 2.9000 1.3400 2.9000 1.1000 3.0200 1.1000 3.0200 1.2200 3.6200 1.2200 ;
        POLYGON  3.5000 2.2100 3.3800 2.2100 3.3800 1.5800 2.7800 1.5800 2.7800 1.6200 1.5100 1.6200
                 1.5100 1.3700 1.6300 1.3700 1.6300 1.5000 2.6600 1.5000 2.6600 0.7200 2.6300 0.7200
                 2.6300 0.6000 2.8700 0.6000 2.8700 0.7200 2.7800 0.7200 2.7800 1.4600 3.5000 1.4600 ;
        POLYGON  3.0800 2.2100 2.9600 2.2100 2.9600 1.8600 2.1900 1.8600 2.1900 2.2100 2.0700 2.2100
                 2.0700 1.7400 2.9600 1.7400 2.9600 1.7000 3.0800 1.7000 ;
        POLYGON  2.2700 1.1000 1.3500 1.1000 1.3500 2.2100 1.2300 2.2100 1.2300 1.1000 0.8000 1.1000
                 0.8000 1.2200 0.6800 1.2200 0.6800 0.9800 1.2300 0.9800 1.2300 0.5400 1.3500 0.5400
                 1.3500 0.9800 2.1500 0.9800 2.1500 0.8600 2.2700 0.8600 ;
    END
END DFFSHQX1

MACRO DFFRXL
    CLASS CORE ;
    FOREIGN DFFRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 0.9200 7.5250 1.1900 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.2200 2.0150 1.4500 ;
        RECT  1.8150 1.1800 1.9350 1.5900 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3384  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 2.8200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 1.1500 3.2150 1.3800 ;
        RECT  2.9150 1.1500 3.1750 1.4050 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1584  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 0.7000 1.4850 0.8200 ;
        RECT  1.3650 0.5800 1.4850 0.8200 ;
        RECT  1.2150 1.4650 1.3800 1.7250 ;
        RECT  1.2150 0.7000 1.3350 2.0900 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.2650 0.6800 7.5050 0.8000 ;
        RECT  7.3850 -0.1800 7.5050 0.8000 ;
        RECT  5.3750 0.4700 5.6150 0.5900 ;
        RECT  5.4950 -0.1800 5.6150 0.5900 ;
        RECT  3.3150 -0.1800 3.4350 0.7500 ;
        RECT  1.7850 -0.1800 1.9050 0.8200 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.6650 2.1100 7.7850 2.7900 ;
        RECT  6.0650 2.1500 6.1850 2.7900 ;
        RECT  5.2550 2.2900 5.4950 2.7900 ;
        RECT  3.3150 2.2900 3.5550 2.7900 ;
        RECT  2.4450 2.1500 2.5650 2.7900 ;
        RECT  1.6950 2.2300 1.8150 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.3250 1.7500 8.0850 1.7500 8.0850 1.4300 7.2250 1.4300 7.2250 1.5500 7.1050 1.5500
                 7.1050 1.4300 7.0250 1.4300 7.0250 0.5000 5.8550 0.5000 5.8550 0.8300 5.1350 0.8300
                 5.1350 0.4800 4.6550 0.4800 4.6550 1.0600 3.9950 1.0600 3.9950 1.4100 3.8750 1.4100
                 3.8750 0.9400 4.5350 0.9400 4.5350 0.3600 5.2550 0.3600 5.2550 0.7100 5.7350 0.7100
                 5.7350 0.3800 6.2350 0.3800 6.2350 0.3600 6.4750 0.3600 6.4750 0.3800 7.1450 0.3800
                 7.1450 1.3100 7.8250 1.3100 7.8250 0.6200 7.9450 0.6200 7.9450 1.3100 8.2050 1.3100
                 8.2050 1.6300 8.3250 1.6300 ;
        POLYGON  8.1250 2.2500 8.0050 2.2500 8.0050 1.9900 7.3300 1.9900 7.3300 2.1500 6.9200 2.1500
                 6.9200 2.2500 6.6800 2.2500 6.6800 2.1500 6.3050 2.1500 6.3050 2.0300 5.9350 2.0300
                 5.9350 1.9300 2.1750 1.9300 2.1750 1.9500 2.0550 1.9500 2.0550 1.7100 2.2650 1.7100
                 2.2650 0.6000 2.3850 0.6000 2.3850 1.8100 4.5350 1.8100 4.5350 1.3300 4.7550 1.3300
                 4.7550 1.1900 4.8750 1.1900 4.8750 1.4500 4.6550 1.4500 4.6550 1.8100 6.0550 1.8100
                 6.0550 1.9100 6.4250 1.9100 6.4250 2.0300 7.2100 2.0300 7.2100 1.8700 8.1250 1.8700 ;
        POLYGON  7.0850 1.9100 6.9650 1.9100 6.9650 1.7900 6.7850 1.7900 6.7850 1.3700 5.2350 1.3700
                 5.2350 1.2500 6.5450 1.2500 6.5450 0.6200 6.6650 0.6200 6.6650 1.2500 6.9050 1.2500
                 6.9050 1.6700 7.0850 1.6700 ;
        POLYGON  6.6650 1.8700 6.5450 1.8700 6.5450 1.6900 5.7350 1.6900 5.7350 1.5700 6.6650 1.5700 ;
        POLYGON  6.2250 1.1300 5.1150 1.1300 5.1150 1.6900 4.7750 1.6900 4.7750 1.5700 4.9950 1.5700
                 4.9950 1.0700 4.7750 1.0700 4.7750 0.6000 5.0150 0.6000 5.0150 0.9500 5.1150 0.9500
                 5.1150 1.0100 6.2250 1.0100 ;
        RECT  2.9950 2.0500 5.8150 2.1700 ;
        POLYGON  4.4150 0.7200 3.7550 0.7200 3.7550 1.5300 4.0950 1.5300 4.0950 1.5700 4.2150 1.5700
                 4.2150 1.6900 3.9750 1.6900 3.9750 1.6500 3.6350 1.6500 3.6350 1.0300 2.7450 1.0300
                 2.7450 0.9100 3.6350 0.9100 3.6350 0.6000 4.4150 0.6000 ;
        POLYGON  3.5150 1.6450 3.0750 1.6450 3.0750 1.6900 2.8350 1.6900 2.8350 1.6450 2.5050 1.6450
                 2.5050 0.6300 2.6750 0.6300 2.6750 0.4800 2.1450 0.4800 2.1450 1.0600 1.6950 1.0600
                 1.6950 1.1000 1.4550 1.1000 1.4550 0.9400 2.0250 0.9400 2.0250 0.3600 2.7950 0.3600
                 2.7950 0.7500 2.6250 0.7500 2.6250 1.5250 3.3950 1.5250 3.3950 1.1900 3.5150 1.1900 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFRXL

MACRO DFFRX4
    CLASS CORE ;
    FOREIGN DFFRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.4300 0.4050 1.5500 ;
        RECT  0.2850 1.1250 0.4050 1.5500 ;
        RECT  0.0700 1.4300 0.2200 1.8400 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.0200 1.6650 1.1400 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        RECT  1.2600 1.0200 1.3800 1.4350 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5350 0.9300 6.6950 1.0500 ;
        RECT  5.5350 0.6300 5.6550 1.0900 ;
        RECT  5.0350 0.6300 5.6550 0.7500 ;
        RECT  5.0350 0.3800 5.1550 0.7500 ;
        RECT  3.9550 0.3800 5.1550 0.5000 ;
        RECT  3.0850 1.2400 4.0750 1.3600 ;
        RECT  3.9550 0.3800 4.0750 1.3600 ;
        RECT  3.9250 0.9400 4.0750 1.3600 ;
        RECT  3.7850 0.9400 4.0750 1.0900 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.1550 0.6800 8.3550 0.8000 ;
        RECT  8.1750 1.3200 8.2950 2.2100 ;
        RECT  7.3200 1.3200 8.2950 1.4400 ;
        RECT  7.3200 1.1750 7.4700 1.4400 ;
        RECT  7.3200 0.6800 7.4400 1.5600 ;
        RECT  7.2150 1.4400 7.3350 2.2100 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0750 0.6800 10.2750 0.8000 ;
        RECT  9.8950 1.5400 10.0150 2.2100 ;
        RECT  9.8550 1.3200 9.9750 1.6600 ;
        RECT  9.0600 1.3200 9.9750 1.4400 ;
        RECT  9.0900 0.6800 9.2100 1.5600 ;
        RECT  9.0550 1.4400 9.1750 2.2100 ;
        RECT  9.0600 1.1750 9.2100 1.5600 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.6350 -0.1800 10.7550 0.6700 ;
        RECT  9.5550 -0.1800 9.7950 0.3200 ;
        RECT  8.5950 -0.1800 8.8350 0.3200 ;
        RECT  7.6350 -0.1800 7.8750 0.3200 ;
        RECT  6.6750 -0.1800 6.9150 0.3200 ;
        RECT  5.2750 0.3900 5.5150 0.5100 ;
        RECT  5.3950 -0.1800 5.5150 0.5100 ;
        RECT  3.5950 0.6800 3.8350 0.8000 ;
        RECT  3.7150 -0.1800 3.8350 0.8000 ;
        RECT  1.6850 0.5400 1.9250 0.6600 ;
        RECT  1.6850 -0.1800 1.8050 0.6600 ;
        RECT  1.2950 0.5400 1.5350 0.6600 ;
        RECT  1.2950 -0.1800 1.4150 0.6600 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.3150 1.5600 10.4350 2.7900 ;
        RECT  9.4750 1.5600 9.5950 2.7900 ;
        RECT  8.6350 1.5600 8.7550 2.7900 ;
        RECT  7.7550 1.5600 7.8750 2.7900 ;
        RECT  6.7950 1.7300 6.9150 2.7900 ;
        RECT  5.9550 1.7300 6.0750 2.7900 ;
        RECT  5.1150 1.7300 5.2350 2.7900 ;
        RECT  3.7350 2.2900 3.9750 2.7900 ;
        RECT  2.5350 2.2000 2.7750 2.7900 ;
        RECT  1.2850 2.2300 1.4050 2.7900 ;
        RECT  0.1350 1.9700 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.1750 0.8600 10.9950 0.8600 10.9950 1.4200 10.8550 1.4200 10.8550 2.2100
                 10.7350 2.2100 10.7350 1.4200 10.0950 1.4200 10.0950 1.2800 10.3350 1.2800
                 10.3350 1.3000 10.8750 1.3000 10.8750 0.7400 11.0550 0.7400 11.0550 0.6200
                 11.1750 0.6200 ;
        POLYGON  10.7150 1.1800 10.5950 1.1800 10.5950 0.9100 10.3950 0.9100 10.3950 0.5600
                 8.5950 0.5600 8.5950 1.0800 8.5550 1.0800 8.5550 1.2000 8.4350 1.2000 8.4350 0.9600
                 8.4750 0.9600 8.4750 0.5600 6.2150 0.5600 6.2150 0.6100 5.9750 0.6100 5.9750 0.4900
                 6.0950 0.4900 6.0950 0.4400 10.5150 0.4400 10.5150 0.7900 10.7150 0.7900 ;
        POLYGON  7.0550 1.6100 6.4950 1.6100 6.4950 2.2100 6.3750 2.2100 6.3750 1.6100 5.6550 1.6100
                 5.6550 2.2100 5.5350 2.2100 5.5350 1.6100 5.0550 1.6100 5.0550 1.5500 4.9350 1.5500
                 4.9350 1.4300 5.1750 1.4300 5.1750 1.4900 6.9350 1.4900 6.9350 1.2400 7.0550 1.2400 ;
        POLYGON  5.9150 1.3700 5.2950 1.3700 5.2950 0.9900 4.5750 0.9900 4.5750 1.9700 4.4550 1.9700
                 4.4550 0.7500 4.6150 0.7500 4.6150 0.6200 4.7350 0.6200 4.7350 0.8700 5.4150 0.8700
                 5.4150 1.2500 5.9150 1.2500 ;
        POLYGON  4.9350 1.2300 4.8150 1.2300 4.8150 2.2100 4.3750 2.2100 4.3750 2.2300 4.1350 2.2300
                 4.1350 2.2100 4.0950 2.2100 4.0950 2.1700 3.6150 2.1700 3.6150 2.2500 2.8950 2.2500
                 2.8950 2.0800 2.3900 2.0800 2.3900 2.2200 2.1500 2.2200 2.1500 2.1100 1.0650 2.1100
                 1.0650 2.2500 0.9450 2.2500 0.9450 2.1100 0.6750 2.1100 0.6750 2.2000 0.5550 2.2000
                 0.5550 2.0800 0.5450 2.0800 0.5450 0.6800 0.6650 0.6800 0.6650 1.9600 0.6750 1.9600
                 0.6750 1.9900 2.0050 1.9900 2.0050 1.9600 3.0150 1.9600 3.0150 2.1300 3.4950 2.1300
                 3.4950 2.0500 4.2150 2.0500 4.2150 2.0900 4.6950 2.0900 4.6950 1.1100 4.9350 1.1100 ;
        POLYGON  4.3150 1.7200 4.1550 1.7200 4.1550 1.8500 4.0350 1.8500 4.0350 1.6000 2.7650 1.6000
                 2.7650 1.4800 4.1950 1.4800 4.1950 0.6200 4.3150 0.6200 ;
        POLYGON  3.6650 1.1200 2.5050 1.1200 2.5050 1.4800 2.2850 1.4800 2.2850 1.7000 2.1050 1.7000
                 2.1050 1.8400 1.9850 1.8400 1.9850 1.5800 2.1650 1.5800 2.1650 1.3600 2.3850 1.3600
                 2.3850 0.6800 2.6250 0.6800 2.6250 0.8000 2.5050 0.8000 2.5050 1.0000 3.6650 1.0000 ;
        POLYGON  3.5950 0.4800 2.1650 0.4800 2.1650 0.9000 1.9050 0.9000 1.9050 1.3400 2.0250 1.3400
                 2.0250 1.4600 1.7850 1.4600 1.7850 0.9000 1.0550 0.9000 1.0550 1.6900 0.9850 1.6900
                 0.9850 1.8100 0.8650 1.8100 0.8650 1.5700 0.9350 1.5700 0.9350 0.4800 1.0550 0.4800
                 1.0550 0.7800 2.0450 0.7800 2.0450 0.3600 3.5950 0.3600 ;
        POLYGON  3.3750 2.0100 3.1350 2.0100 3.1350 1.8400 2.4050 1.8400 2.4050 1.6000 2.5250 1.6000
                 2.5250 1.7200 3.2550 1.7200 3.2550 1.8900 3.3750 1.8900 ;
    END
END DFFRX4

MACRO DFFRX2
    CLASS CORE ;
    FOREIGN DFFRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.4500 0.8550 1.6800 ;
        RECT  0.7150 1.1600 0.8350 1.6800 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4750 1.2700 2.7150 1.4400 ;
        RECT  2.3350 1.2300 2.5950 1.4300 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.8150 1.4500 6.0750 1.6700 ;
        RECT  5.8250 1.2800 5.9450 1.6700 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7150 1.4650 6.8900 1.7250 ;
        RECT  6.7150 0.8000 6.8350 2.1500 ;
        RECT  6.5250 0.8000 6.8350 0.9200 ;
        RECT  6.5250 0.6800 6.6450 0.9200 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5550 1.4650 7.7600 1.7250 ;
        RECT  7.5550 1.4650 7.6750 2.1500 ;
        RECT  7.4250 0.7400 7.6650 0.8600 ;
        RECT  7.4650 0.7400 7.5850 1.6200 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  7.9050 -0.1800 8.1450 0.3200 ;
        RECT  6.9450 -0.1800 7.1850 0.3200 ;
        RECT  6.0450 -0.1800 6.1650 0.9200 ;
        RECT  4.2250 -0.1800 4.3450 0.8600 ;
        RECT  2.5050 0.5100 2.7450 0.6300 ;
        RECT  2.5050 -0.1800 2.6250 0.6300 ;
        RECT  0.9450 0.6800 1.1850 0.8000 ;
        RECT  0.9450 -0.1800 1.0650 0.8000 ;
        RECT  0.5550 -0.1800 0.6750 0.8000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  7.9750 1.5000 8.0950 2.7900 ;
        RECT  7.1350 1.5000 7.2550 2.7900 ;
        RECT  6.2950 1.7900 6.4150 2.7900 ;
        RECT  5.4850 2.0800 5.6050 2.7900 ;
        RECT  4.5250 2.0800 4.6450 2.7900 ;
        RECT  2.9250 2.0400 3.0450 2.7900 ;
        RECT  1.8450 2.2900 2.0850 2.7900 ;
        RECT  0.6150 2.1200 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.5650 1.3450 8.5150 1.3450 8.5150 1.7400 8.3950 1.7400 8.3950 1.3450 7.7050 1.3450
                 7.7050 1.2250 8.4450 1.2250 8.4450 0.6800 8.5650 0.6800 ;
        POLYGON  8.5050 0.5200 8.3850 0.5200 8.3850 0.5600 7.0750 0.5600 7.0750 1.2600 6.9550 1.2600
                 6.9550 0.5600 6.4050 0.5600 6.4050 1.2400 6.2850 1.2400 6.2850 1.1600 5.8050 1.1600
                 5.8050 0.5600 5.2850 0.5600 5.2850 0.6800 5.4450 0.6800 5.4450 1.3600 5.1250 1.3600
                 5.1250 1.7200 5.0050 1.7200 5.0050 1.3600 4.5050 1.3600 4.5050 1.3400 4.3850 1.3400
                 4.3850 1.2200 4.6250 1.2200 4.6250 1.2400 5.3250 1.2400 5.3250 0.8000 5.1650 0.8000
                 5.1650 0.4400 5.9250 0.4400 5.9250 1.0400 6.2850 1.0400 6.2850 0.4400 8.2650 0.4400
                 8.2650 0.4000 8.5050 0.4000 ;
        POLYGON  5.9950 2.0300 5.8750 2.0300 5.8750 1.9600 4.4050 1.9600 4.4050 2.2300 3.8650 2.2300
                 3.8650 2.2500 3.6250 2.2500 3.6250 2.2300 3.1650 2.2300 3.1650 1.9200 2.8050 1.9200
                 2.8050 2.1700 1.3850 2.1700 1.3850 2.1000 0.8550 2.1000 0.8550 2.0000 0.3950 2.0000
                 0.3950 2.1600 0.2750 2.1600 0.2750 1.8800 0.9750 1.8800 0.9750 1.9800 1.6250 1.9800
                 1.6250 2.0500 2.6850 2.0500 2.6850 1.8000 3.2850 1.8000 3.2850 2.1100 4.2850 2.1100
                 4.2850 1.8400 5.5650 1.8400 5.5650 0.6800 5.6850 0.6800 5.6850 1.7900 5.9950 1.7900 ;
        POLYGON  5.2050 1.1200 4.9650 1.1200 4.9650 1.1000 4.2650 1.1000 4.2650 1.7200 4.0050 1.7200
                 4.0050 1.8100 3.7650 1.8100 3.7650 1.6900 3.8850 1.6900 3.8850 1.6000 4.1450 1.6000
                 4.1450 1.1000 3.5850 1.1000 3.5850 0.6200 3.7050 0.6200 3.7050 0.9800 5.0850 0.9800
                 5.0850 1.0000 5.2050 1.0000 ;
        POLYGON  4.0250 1.4800 3.9050 1.4800 3.9050 1.3600 3.3450 1.3600 3.3450 0.5000 2.9850 0.5000
                 2.9850 0.8700 2.2650 0.8700 2.2650 0.5600 1.4250 0.5600 1.4250 1.0400 1.1950 1.0400
                 1.1950 1.4000 1.0750 1.4000 1.0750 1.0400 0.2550 1.0400 0.2550 1.7200 0.1350 1.7200
                 0.1350 0.7400 0.0750 0.7400 0.0750 0.6200 0.3150 0.6200 0.3150 0.7400 0.2550 0.7400
                 0.2550 0.9200 1.3050 0.9200 1.3050 0.4400 1.7250 0.4400 1.7250 0.3600 1.9650 0.3600
                 1.9650 0.4400 2.3850 0.4400 2.3850 0.7500 2.8650 0.7500 2.8650 0.3800 3.4650 0.3800
                 3.4650 1.2400 4.0250 1.2400 ;
        POLYGON  3.5250 1.9900 3.4050 1.9900 3.4050 1.6800 2.0950 1.6800 2.0950 1.4100 2.2150 1.4100
                 2.2150 1.5600 3.1050 1.5600 3.1050 0.6200 3.2250 0.6200 3.2250 1.5600 3.5250 1.5600 ;
        POLYGON  2.9850 1.1200 2.7150 1.1200 2.7150 1.1100 1.7050 1.1100 1.7050 1.4800 1.5150 1.4800
                 1.5150 1.6400 1.3350 1.6400 1.3350 1.7600 1.2150 1.7600 1.2150 1.5200 1.3950 1.5200
                 1.3950 1.3600 1.5850 1.3600 1.5850 0.6800 1.8250 0.6800 1.8250 0.8000 1.7050 0.8000
                 1.7050 0.9900 2.8350 0.9900 2.8350 1.0000 2.9850 1.0000 ;
        POLYGON  2.5650 1.9300 2.0600 1.9300 2.0600 1.9200 1.7950 1.9200 1.7950 1.8600 1.6350 1.8600
                 1.6350 1.6000 1.7550 1.6000 1.7550 1.7400 1.9150 1.7400 1.9150 1.8000 2.1800 1.8000
                 2.1800 1.8100 2.5650 1.8100 ;
    END
END DFFRX2

MACRO DFFRX1
    CLASS CORE ;
    FOREIGN DFFRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2650 0.9200 7.5250 1.1900 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.2550 2.1050 1.4600 ;
        RECT  1.7550 1.2300 2.0150 1.4600 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.3312  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 2.7600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 1.1950 3.2750 1.3950 ;
        RECT  2.9150 1.1700 3.1750 1.3950 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2888  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3750 0.6100 1.4950 0.8700 ;
        RECT  1.2850 1.2300 1.4050 2.2100 ;
        RECT  1.2650 0.7500 1.3850 1.3500 ;
        RECT  1.2300 0.8850 1.3850 1.1450 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.2650 0.6800 7.5050 0.8000 ;
        RECT  7.3850 -0.1800 7.5050 0.8000 ;
        RECT  5.4250 0.4700 5.6650 0.5900 ;
        RECT  5.5450 -0.1800 5.6650 0.5900 ;
        RECT  3.3150 0.6100 3.5550 0.7300 ;
        RECT  3.4350 -0.1800 3.5550 0.7300 ;
        RECT  1.7350 0.6700 1.9750 0.7900 ;
        RECT  1.7350 -0.1800 1.8550 0.7900 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.6650 2.1100 7.7850 2.7900 ;
        RECT  6.0650 2.1500 6.1850 2.7900 ;
        RECT  5.2550 2.2900 5.4950 2.7900 ;
        RECT  3.3750 2.2900 3.6150 2.7900 ;
        RECT  2.5150 2.1500 2.6350 2.7900 ;
        RECT  1.7650 2.2000 1.8850 2.7900 ;
        RECT  0.6150 1.9800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.3250 1.7500 8.0850 1.7500 8.0850 1.4300 7.2250 1.4300 7.2250 1.5500 7.1050 1.5500
                 7.1050 1.4300 7.0250 1.4300 7.0250 0.5000 5.9050 0.5000 5.9050 0.8300 5.1850 0.8300
                 5.1850 0.4900 4.7050 0.4900 4.7050 1.0700 4.0550 1.0700 4.0550 1.4100 3.9350 1.4100
                 3.9350 0.9500 4.5850 0.9500 4.5850 0.3700 5.3050 0.3700 5.3050 0.7100 5.7850 0.7100
                 5.7850 0.3800 6.2350 0.3800 6.2350 0.3600 6.4750 0.3600 6.4750 0.3800 7.1450 0.3800
                 7.1450 1.3100 7.8250 1.3100 7.8250 0.6200 7.9450 0.6200 7.9450 1.3100 8.2050 1.3100
                 8.2050 1.6300 8.3250 1.6300 ;
        POLYGON  8.1250 2.2500 8.0050 2.2500 8.0050 1.9900 7.3300 1.9900 7.3300 2.1500 6.9200 2.1500
                 6.9200 2.2500 6.6800 2.2500 6.6800 2.1500 6.3050 2.1500 6.3050 1.9300 2.1250 1.9300
                 2.1250 1.5800 2.3350 1.5800 2.3350 0.6100 2.4550 0.6100 2.4550 1.8100 4.5950 1.8100
                 4.5950 1.3100 4.8150 1.3100 4.8150 1.1900 4.9350 1.1900 4.9350 1.4300 4.7150 1.4300
                 4.7150 1.8100 6.4250 1.8100 6.4250 2.0300 7.2100 2.0300 7.2100 1.8700 8.1250 1.8700 ;
        POLYGON  7.0850 1.9100 6.9650 1.9100 6.9650 1.7900 6.8650 1.7900 6.8650 1.6700 6.7850 1.6700
                 6.7850 1.3600 5.4150 1.3600 5.4150 1.4300 5.2950 1.4300 5.2950 1.1900 5.4150 1.1900
                 5.4150 1.2400 6.5450 1.2400 6.5450 0.6200 6.6650 0.6200 6.6650 1.2400 6.9050 1.2400
                 6.9050 1.5500 6.9850 1.5500 6.9850 1.6700 7.0850 1.6700 ;
        POLYGON  6.6650 1.8700 6.5450 1.8700 6.5450 1.6900 5.7350 1.6900 5.7350 1.5700 6.6650 1.5700 ;
        POLYGON  6.2250 1.1200 5.9850 1.1200 5.9850 1.0700 5.1750 1.0700 5.1750 1.6900 4.8350 1.6900
                 4.8350 1.5700 5.0550 1.5700 5.0550 1.0700 4.8250 1.0700 4.8250 0.6100 5.0650 0.6100
                 5.0650 0.9500 6.1050 0.9500 6.1050 1.0000 6.2250 1.0000 ;
        RECT  3.0550 2.0500 5.8150 2.1700 ;
        POLYGON  4.4650 0.7300 3.8150 0.7300 3.8150 1.5300 4.1550 1.5300 4.1550 1.5700 4.2750 1.5700
                 4.2750 1.6900 4.0350 1.6900 4.0350 1.6500 3.6950 1.6500 3.6950 1.0500 2.8150 1.0500
                 2.8150 0.9300 3.6950 0.9300 3.6950 0.6100 4.4650 0.6100 ;
        POLYGON  3.5750 1.6350 3.1350 1.6350 3.1350 1.6900 2.8950 1.6900 2.8950 1.6350 2.5750 1.6350
                 2.5750 0.6700 2.7350 0.6700 2.7350 0.4900 2.2150 0.4900 2.2150 1.1100 1.5050 1.1100
                 1.5050 0.9900 2.0950 0.9900 2.0950 0.3700 2.8550 0.3700 2.8550 0.7900 2.6950 0.7900
                 2.6950 1.5150 3.4550 1.5150 3.4550 1.1900 3.5750 1.1900 ;
        POLYGON  1.1050 0.9200 1.0950 0.9200 1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000
                 0.3750 1.0800 0.9750 1.0800 0.9750 0.8000 0.9850 0.8000 0.9850 0.6800 1.1050 0.6800 ;
    END
END DFFRX1

MACRO DFFRHQX8
    CLASS CORE ;
    FOREIGN DFFRHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.1800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6450 0.7250 2.9650 0.8450 ;
        RECT  2.6650 1.3400 2.7850 2.0850 ;
        RECT  2.6450 0.7250 2.7650 1.4600 ;
        RECT  0.2650 1.0250 2.7650 1.1450 ;
        RECT  1.9450 0.6650 2.0650 1.4600 ;
        RECT  1.8250 1.3400 1.9450 2.0850 ;
        RECT  1.1050 0.6650 1.2250 1.4600 ;
        RECT  0.9850 1.3400 1.1050 2.0800 ;
        RECT  0.2650 0.8850 0.5100 1.1450 ;
        RECT  0.2650 0.6650 0.3850 1.4600 ;
        RECT  0.1450 1.3400 0.2650 2.0800 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.8850 0.8600 11.1250 1.0400 ;
        RECT  10.7450 0.8850 11.0050 1.0900 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.4140  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4100  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.0098  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.5850 0.3600 4.7050 1.1600 ;
        RECT  3.4450 0.3600 4.7050 0.4800 ;
        RECT  3.4450 0.3600 3.5650 1.1800 ;
        RECT  3.2600 0.8850 3.5650 1.1450 ;
        END
    END RN
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.6150 1.1100 11.8750 1.3800 ;
        RECT  11.5750 1.1100 11.8750 1.3600 ;
        END
    END CK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 12.1800 0.1800 ;
        RECT  11.3750 -0.1800 11.4950 0.7500 ;
        RECT  10.9250 0.5000 11.1650 0.6200 ;
        RECT  10.9250 -0.1800 11.0450 0.6200 ;
        RECT  8.7750 0.4300 9.0150 0.5500 ;
        RECT  8.8950 -0.1800 9.0150 0.5500 ;
        RECT  6.3950 -0.1800 6.6350 0.3200 ;
        RECT  4.8250 -0.1800 4.9450 0.6500 ;
        RECT  3.2050 -0.1800 3.3250 0.6500 ;
        RECT  2.3650 -0.1800 2.4850 0.6550 ;
        RECT  1.5250 -0.1800 1.6450 0.6550 ;
        RECT  0.6850 -0.1800 0.8050 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 12.1800 2.7900 ;
        RECT  11.1850 1.7400 11.3050 2.7900 ;
        RECT  9.6750 2.2900 9.9150 2.7900 ;
        RECT  8.7750 2.0100 8.8950 2.7900 ;
        RECT  8.6550 2.0100 8.8950 2.1300 ;
        RECT  6.6350 2.2200 6.8750 2.7900 ;
        RECT  5.7850 2.2200 6.0250 2.7900 ;
        RECT  4.8250 1.9000 5.0650 2.0200 ;
        RECT  4.8250 1.9000 4.9450 2.7900 ;
        RECT  3.8650 1.9000 4.1050 2.0200 ;
        RECT  3.8650 1.9000 3.9850 2.7900 ;
        RECT  3.0850 1.5400 3.2050 2.7900 ;
        RECT  2.2450 1.3400 2.3650 2.7900 ;
        RECT  1.4050 1.3400 1.5250 2.7900 ;
        RECT  0.5650 1.3400 0.6850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.9150 0.9900 11.4550 0.9900 11.4550 1.5000 11.5450 1.5000 11.5450 1.6400
                 11.7250 1.6400 11.7250 1.8800 11.6050 1.8800 11.6050 1.7600 11.4250 1.7600
                 11.4250 1.6200 11.3350 1.6200 11.3350 1.3600 10.2650 1.3600 10.2650 1.3100
                 10.1250 1.3100 10.1250 1.1900 10.3850 1.1900 10.3850 1.2400 11.3350 1.2400
                 11.3350 0.8700 11.7950 0.8700 11.7950 0.5100 11.9150 0.5100 ;
        POLYGON  10.6650 1.9900 10.5450 1.9900 10.5450 1.6000 9.8850 1.6000 9.8850 1.5600 8.6950 1.5600
                 8.6950 1.1500 8.8150 1.1500 8.8150 1.4400 9.8850 1.4400 9.8850 0.6000 10.1250 0.6000
                 10.1250 0.7200 10.0050 0.7200 10.0050 1.4800 10.6650 1.4800 ;
        POLYGON  10.6250 1.1200 10.5050 1.1200 10.5050 0.4800 9.7650 0.4800 9.7650 1.1000 9.6450 1.1000
                 9.6450 0.7400 9.5000 0.7400 9.5000 0.7900 8.5350 0.7900 8.5350 0.4800 7.9550 0.4800
                 7.9550 0.9200 7.9750 0.9200 7.9750 1.0400 7.7350 1.0400 7.7350 0.9200 7.8350 0.9200
                 7.8350 0.4800 7.3550 0.4800 7.3550 1.5400 6.3750 1.5400 6.3750 1.6200 6.0350 1.6200
                 6.0350 0.8000 5.9150 0.8000 5.9150 0.6800 6.1550 0.6800 6.1550 1.4200 7.2350 1.4200
                 7.2350 0.3600 8.6550 0.3600 8.6550 0.6700 9.3800 0.6700 9.3800 0.6200 9.6450 0.6200
                 9.6450 0.3600 10.6250 0.3600 ;
        POLYGON  10.4450 2.2500 10.2050 2.2500 10.2050 2.1700 9.0150 2.1700 9.0150 1.8900 7.9350 1.8900
                 7.9350 1.2100 8.3350 1.2100 8.3350 1.3300 8.0550 1.3300 8.0550 1.7700 9.1350 1.7700
                 9.1350 2.0500 10.3250 2.0500 10.3250 2.1300 10.4450 2.1300 ;
        POLYGON  10.3050 1.9300 9.2550 1.9300 9.2550 1.6900 9.3750 1.6900 9.3750 1.8100 10.0650 1.8100
                 10.0650 1.7200 10.3050 1.7200 ;
        POLYGON  9.4050 1.3200 9.2850 1.3200 9.2850 1.0300 8.5750 1.0300 8.5750 1.6500 8.1750 1.6500
                 8.1750 1.5300 8.4550 1.5300 8.4550 1.0300 8.1750 1.0300 8.1750 0.6000 8.4150 0.6000
                 8.4150 0.9100 9.4050 0.9100 ;
        POLYGON  8.3350 2.2500 7.8300 2.2500 7.8300 2.2300 7.2350 2.2300 7.2350 2.1000 5.4250 2.1000
                 5.4250 2.2500 5.1850 2.2500 5.1850 2.1300 5.3050 2.1300 5.3050 1.9800 7.3550 1.9800
                 7.3550 2.1100 7.9500 2.1100 7.9500 2.1300 8.3350 2.1300 ;
        POLYGON  7.7150 0.7200 7.5950 0.7200 7.5950 1.9900 7.4750 1.9900 7.4750 1.8600 5.6650 1.8600
                 5.6650 1.7800 4.0650 1.7800 4.0650 1.0400 4.1850 1.0400 4.1850 1.6600 5.6650 1.6600
                 5.6650 1.2600 5.6450 1.2600 5.6450 1.0200 5.7850 1.0200 5.7850 1.7400 7.4750 1.7400
                 7.4750 0.6000 7.7150 0.6000 ;
        POLYGON  7.1150 1.3000 6.2750 1.3000 6.2750 1.1800 6.9950 1.1800 6.9950 0.8800 7.1150 0.8800 ;
        POLYGON  6.8550 1.0600 6.6150 1.0600 6.6150 0.5600 5.7050 0.5600 5.7050 0.9000 5.4250 0.9000
                 5.4250 1.4000 5.5450 1.4000 5.5450 1.5400 5.3050 1.5400 5.3050 1.4000 4.5850 1.4000
                 4.5850 1.5400 4.3450 1.5400 4.3450 0.9200 3.9450 0.9200 3.9450 1.4200 3.6250 1.4200
                 3.6250 2.0800 3.5050 2.0800 3.5050 1.4200 3.0200 1.4200 3.0200 1.2000 2.8850 1.2000
                 2.8850 1.0800 3.1400 1.0800 3.1400 1.3000 3.8250 1.3000 3.8250 0.7200 3.9250 0.7200
                 3.9250 0.6000 4.0450 0.6000 4.0450 0.8000 4.4650 0.8000 4.4650 1.2800 5.3050 1.2800
                 5.3050 0.7800 5.5850 0.7800 5.5850 0.4400 6.7350 0.4400 6.7350 0.9400 6.8550 0.9400 ;
    END
END DFFRHQX8

MACRO DFFRHQX4
    CLASS CORE ;
    FOREIGN DFFRHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9350 1.4900 2.1750 1.6100 ;
        RECT  1.9350 1.3150 2.1400 1.6100 ;
        RECT  2.0200 0.6300 2.1400 1.6100 ;
        RECT  1.2300 1.3150 2.1400 1.4350 ;
        RECT  1.1800 1.1750 1.3800 1.3150 ;
        RECT  0.9750 1.4900 1.3500 1.6100 ;
        RECT  1.2300 1.1750 1.3500 1.6100 ;
        RECT  1.1800 0.6300 1.3000 1.3150 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.8800 0.9300 9.0000 1.2400 ;
        RECT  8.7700 0.8300 8.9200 1.1450 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.1100 0.8550 1.3800 ;
        RECT  0.4950 1.1100 0.8550 1.3600 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2580  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7550 1.1600 6.5350 1.2800 ;
        RECT  6.4150 1.0400 6.5350 1.2800 ;
        RECT  5.7550 0.3600 5.8750 1.2800 ;
        RECT  4.6150 0.3600 5.8750 0.4800 ;
        RECT  3.5050 0.7300 4.7350 0.8500 ;
        RECT  4.6150 0.3600 4.7350 0.8500 ;
        RECT  3.6950 0.7300 3.8150 1.1000 ;
        RECT  3.5050 0.3600 3.6250 0.8500 ;
        RECT  2.7100 0.3600 3.6250 0.4800 ;
        RECT  2.7100 0.3600 2.8300 1.1200 ;
        RECT  2.6800 0.5950 2.8300 0.8550 ;
        END
    END RN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  8.9400 -0.1800 9.0600 0.7100 ;
        RECT  5.9950 -0.1800 6.1150 0.6800 ;
        RECT  3.8350 0.4900 4.0750 0.6100 ;
        RECT  3.8350 -0.1800 3.9550 0.6100 ;
        RECT  2.4400 -0.1800 2.5600 0.6800 ;
        RECT  1.6000 -0.1800 1.7200 0.6800 ;
        RECT  0.7600 -0.1800 0.8800 0.8700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  9.0400 1.6000 9.1600 2.7900 ;
        RECT  7.3600 2.2900 7.6000 2.7900 ;
        RECT  5.8600 2.2500 6.1000 2.7900 ;
        RECT  4.2150 1.9400 4.3350 2.7900 ;
        RECT  3.3150 2.2300 3.4350 2.7900 ;
        RECT  2.4750 2.2300 2.5950 2.7900 ;
        RECT  1.4550 1.9700 1.6950 2.0900 ;
        RECT  1.4550 1.9700 1.5750 2.7900 ;
        RECT  0.4950 1.9700 0.7350 2.0900 ;
        RECT  0.4950 1.9700 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.5800 1.8400 9.4600 1.8400 9.4600 1.7200 9.3600 1.7200 9.3600 1.4800 8.7600 1.4800
                 8.7600 2.2000 8.0500 2.2000 8.0500 1.9300 6.6550 1.9300 6.6550 1.8900 5.0950 1.8900
                 5.0950 1.3300 4.6550 1.3300 4.6550 1.2100 5.0950 1.2100 5.0950 1.0000 5.2750 1.0000
                 5.2750 0.8800 5.3950 0.8800 5.3950 1.1200 5.2150 1.1200 5.2150 1.7700 6.7750 1.7700
                 6.7750 1.8100 8.0500 1.8100 8.0500 1.3200 7.6350 1.3200 7.6350 1.1600 7.5150 1.1600
                 7.5150 1.0400 7.7550 1.0400 7.7550 1.2000 8.1700 1.2000 8.1700 2.0800 8.6400 2.0800
                 8.6400 1.3850 8.5300 1.3850 8.5300 1.1000 8.6500 1.1000 8.6500 1.2650 8.7600 1.2650
                 8.7600 1.3600 9.3600 1.3600 9.3600 0.4700 9.4800 0.4700 9.4800 1.6000 9.5800 1.6000 ;
        POLYGON  8.5200 1.9600 8.4000 1.9600 8.4000 1.6250 8.2900 1.6250 8.2900 0.9200 6.2350 0.9200
                 6.2350 1.0400 5.9950 1.0400 5.9950 0.8000 7.7350 0.8000 7.7350 0.5400 7.8550 0.5400
                 7.8550 0.8000 8.4100 0.8000 8.4100 1.5050 8.5200 1.5050 ;
        POLYGON  7.9300 1.6900 7.8100 1.6900 7.8100 1.6500 7.1350 1.6500 7.1350 1.6900 6.8950 1.6900
                 6.8950 1.5300 7.8100 1.5300 7.8100 1.4400 7.9300 1.4400 ;
        POLYGON  7.9200 2.1700 6.4150 2.1700 6.4150 2.1300 5.7400 2.1300 5.7400 2.2300 5.3150 2.2300
                 5.3150 2.2500 5.0750 2.2500 5.0750 2.2300 4.5600 2.2300 4.5600 1.8200 4.0950 1.8200
                 4.0950 2.1100 1.9900 2.1100 1.9900 1.8500 0.3750 1.8500 0.3750 1.9100 0.2550 1.9100
                 0.2550 2.0300 0.1350 2.0300 0.1350 1.7300 0.2550 1.7300 0.2550 0.6900 0.5200 0.6900
                 0.5200 0.8100 0.3750 0.8100 0.3750 1.7300 2.1100 1.7300 2.1100 1.9900 3.9750 1.9900
                 3.9750 1.7000 4.6800 1.7000 4.6800 2.1100 5.6200 2.1100 5.6200 2.0100 6.5350 2.0100
                 6.5350 2.0500 7.9200 2.0500 ;
        POLYGON  7.3550 1.4100 6.7750 1.4100 6.7750 1.5200 5.6350 1.5200 5.6350 1.6500 5.3350 1.6500
                 5.3350 1.5300 5.5150 1.5300 5.5150 0.7200 5.3750 0.7200 5.3750 0.6000 5.6350 0.6000
                 5.6350 1.4000 6.6550 1.4000 6.6550 1.2900 7.2350 1.2900 7.2350 1.1100 7.3550 1.1100 ;
        POLYGON  5.1950 0.7200 4.9750 0.7200 4.9750 1.0900 4.5350 1.0900 4.5350 1.4500 4.9200 1.4500
                 4.9200 1.5700 4.9750 1.5700 4.9750 1.9900 4.8550 1.9900 4.8550 1.6900 4.8000 1.6900
                 4.8000 1.5700 4.4150 1.5700 4.4150 1.0900 4.0550 1.0900 4.0550 1.3400 3.3350 1.3400
                 3.3350 1.1000 3.4550 1.1000 3.4550 1.2200 3.9350 1.2200 3.9350 0.9700 4.8550 0.9700
                 4.8550 0.6000 5.1950 0.6000 ;
        POLYGON  4.2950 1.5800 3.8550 1.5800 3.8550 1.8700 3.6150 1.8700 3.6150 1.7200 3.7350 1.7200
                 3.7350 1.5800 2.9550 1.5800 2.9550 1.8700 2.8350 1.8700 2.8350 1.3600 2.2750 1.3600
                 2.2750 1.1100 2.3950 1.1100 2.3950 1.2400 2.9550 1.2400 2.9550 1.4600 3.0950 1.4600
                 3.0950 0.6000 3.3750 0.6000 3.3750 0.7200 3.2150 0.7200 3.2150 1.4600 4.1750 1.4600
                 4.1750 1.3400 4.2950 1.3400 ;
    END
END DFFRHQX4

MACRO DFFRHQX2
    CLASS CORE ;
    FOREIGN DFFRHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.1150 0.9000 7.2350 1.3100 ;
        RECT  6.9750 0.9000 7.2350 1.1300 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.1650 1.4750 1.3800 ;
        RECT  1.1850 1.1400 1.4700 1.3800 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 1.2300 3.1750 1.3800 ;
        RECT  2.5950 1.3600 3.0350 1.4800 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6450 1.4650 0.8000 1.7250 ;
        RECT  0.6450 1.4000 0.7700 1.7250 ;
        RECT  0.6450 0.6800 0.7650 2.0500 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.3850 -0.1800 7.5050 0.5400 ;
        RECT  6.8350 0.4200 7.0750 0.5400 ;
        RECT  6.8350 -0.1800 6.9550 0.5400 ;
        RECT  4.9750 0.4300 5.2150 0.5500 ;
        RECT  5.0950 -0.1800 5.2150 0.5500 ;
        RECT  2.6750 0.4600 2.9150 0.5800 ;
        RECT  2.7950 -0.1800 2.9150 0.5800 ;
        RECT  1.0050 0.6600 1.2450 0.7800 ;
        RECT  1.0050 -0.1800 1.1250 0.7800 ;
        RECT  0.2250 -0.1800 0.3450 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.4450 2.2300 7.5650 2.7900 ;
        RECT  5.6550 2.2600 5.8950 2.7900 ;
        RECT  4.5750 2.0100 4.8150 2.1300 ;
        RECT  4.5750 2.0100 4.6950 2.7900 ;
        RECT  2.9750 1.8400 3.0950 2.7900 ;
        RECT  2.8550 1.8400 3.0950 1.9600 ;
        RECT  1.8750 1.7400 1.9950 2.7900 ;
        RECT  1.0650 1.5000 1.1850 2.7900 ;
        RECT  0.2250 1.4000 0.3450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.9850 1.8100 7.8650 1.8100 7.8650 1.5500 6.8250 1.5500 6.8250 1.4300 7.3550 1.4300
                 7.3550 0.7800 6.5600 0.7800 6.5600 0.4800 6.0150 0.4800 6.0150 0.9200 6.1350 0.9200
                 6.1350 1.0400 5.8950 1.0400 5.8950 0.7900 4.7350 0.7900 4.7350 0.4800 4.0950 0.4800
                 4.0950 0.9200 4.3750 0.9200 4.3750 1.0400 3.9750 1.0400 3.9750 0.3600 4.8550 0.3600
                 4.8550 0.6700 5.8950 0.6700 5.8950 0.3600 6.6800 0.3600 6.6800 0.6600 7.4750 0.6600
                 7.4750 1.4300 7.8650 1.4300 7.8650 0.4000 7.9850 0.4000 ;
        POLYGON  7.9050 2.2500 7.7850 2.2500 7.7850 2.1100 7.1100 2.1100 7.1100 2.2500 6.1950 2.2500
                 6.1950 2.1400 4.9350 2.1400 4.9350 1.8900 3.9750 1.8900 3.9750 2.2300 3.2950 2.2300
                 3.2950 1.7200 2.7350 1.7200 2.7350 2.2500 2.1150 2.2500 2.1150 1.6200 1.6050 1.6200
                 1.6050 1.7400 1.4850 1.7400 1.4850 1.5000 1.6050 1.5000 1.6050 0.6000 1.7250 0.6000
                 1.7250 1.5000 2.2350 1.5000 2.2350 2.1300 2.6150 2.1300 2.6150 1.6000 3.2950 1.6000
                 3.2950 1.0600 3.1750 1.0600 3.1750 0.9400 3.4150 0.9400 3.4150 2.1100 3.8550 2.1100
                 3.8550 1.3300 3.7750 1.3300 3.7750 1.2100 4.0150 1.2100 4.0150 1.3300 3.9750 1.3300
                 3.9750 1.7700 5.0550 1.7700 5.0550 2.0200 6.3450 2.0200 6.3450 1.5200 6.2250 1.5200
                 6.2250 1.4000 6.4650 1.4000 6.4650 2.1300 6.9900 2.1300 6.9900 1.9900 7.9050 1.9900 ;
        POLYGON  6.7050 2.0100 6.5850 2.0100 6.5850 1.2800 4.8550 1.2800 4.8550 1.3900 4.7350 1.3900
                 4.7350 1.1500 4.8550 1.1500 4.8550 1.1600 6.2550 1.1600 6.2550 0.7200 6.1350 0.7200
                 6.1350 0.6000 6.3750 0.6000 6.3750 1.1600 6.7050 1.1600 ;
        POLYGON  6.2250 1.9000 6.1050 1.9000 6.1050 1.8700 5.4150 1.8700 5.4150 1.9000 5.1750 1.9000
                 5.1750 1.7500 6.1050 1.7500 6.1050 1.6600 6.2250 1.6600 ;
        POLYGON  5.7750 1.0400 5.5350 1.0400 5.5350 1.0300 4.6150 1.0300 4.6150 1.6500 4.0950 1.6500
                 4.0950 1.5300 4.4950 1.5300 4.4950 0.7200 4.2150 0.7200 4.2150 0.6000 4.6150 0.6000
                 4.6150 0.9100 5.6550 0.9100 5.6550 0.9200 5.7750 0.9200 ;
        POLYGON  3.7350 1.9900 3.6150 1.9900 3.6150 1.5900 3.5350 1.5900 3.5350 0.8200 2.4550 0.8200
                 2.4550 1.0000 2.1750 1.0000 2.1750 0.8800 2.3350 0.8800 2.3350 0.7000 3.5350 0.7000
                 3.5350 0.5000 3.6550 0.5000 3.6550 1.4700 3.7350 1.4700 ;
        POLYGON  3.0550 1.1100 2.6950 1.1100 2.6950 1.2400 2.4750 1.2400 2.4750 2.0100 2.3550 2.0100
                 2.3550 1.2400 1.9350 1.2400 1.9350 0.6000 2.0950 0.6000 2.0950 0.4800 1.4850 0.4800
                 1.4850 1.0200 1.0250 1.0200 1.0250 1.2600 0.9050 1.2600 0.9050 0.9000 1.3650 0.9000
                 1.3650 0.3600 2.2150 0.3600 2.2150 0.7200 2.0550 0.7200 2.0550 1.1200 2.5750 1.1200
                 2.5750 0.9900 3.0550 0.9900 ;
    END
END DFFRHQX2

MACRO DFFRHQX1
    CLASS CORE ;
    FOREIGN DFFRHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5650 0.9600 6.9450 1.2100 ;
        RECT  6.6850 0.9400 6.9450 1.2100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 1.1550 0.9950 1.3200 ;
        RECT  0.5950 1.1850 0.8550 1.3800 ;
        END
    END CK
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1720  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2150 1.2200 2.5950 1.4000 ;
        RECT  2.3350 1.1950 2.5950 1.4000 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 1.3400 0.2550 1.9900 ;
        RECT  0.1350 0.5550 0.2550 0.7950 ;
        RECT  0.0700 1.1750 0.2350 1.4350 ;
        RECT  0.1150 0.6750 0.2350 1.4600 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  7.0350 0.4600 7.2750 0.5800 ;
        RECT  7.0350 -0.1800 7.1550 0.5800 ;
        RECT  6.3550 0.4600 6.5950 0.5800 ;
        RECT  6.3550 -0.1800 6.4750 0.5800 ;
        RECT  4.4950 -0.1800 4.7350 0.3900 ;
        RECT  2.0750 0.4600 2.3150 0.5800 ;
        RECT  2.1950 -0.1800 2.3150 0.5800 ;
        RECT  0.4950 0.6750 0.7350 0.7950 ;
        RECT  0.4950 -0.1800 0.6150 0.7950 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  7.0350 2.1700 7.1550 2.7900 ;
        RECT  5.3750 2.1200 5.4950 2.7900 ;
        RECT  5.2550 2.1200 5.4950 2.2400 ;
        RECT  4.1350 1.7100 4.3750 1.9300 ;
        RECT  4.1350 1.7100 4.2550 2.7900 ;
        RECT  2.5650 1.7600 2.6850 2.7900 ;
        RECT  2.4450 1.7600 2.6850 1.9300 ;
        RECT  1.4350 1.6800 1.5550 2.7900 ;
        RECT  0.5550 1.5000 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.6350 1.8100 7.5150 1.8100 7.5150 1.4500 6.6150 1.4500 6.6150 1.5700 6.4950 1.5700
                 6.4950 1.3300 7.0650 1.3300 7.0650 0.8200 6.1150 0.8200 6.1150 0.4800 5.5350 0.4800
                 5.5350 0.9200 5.6550 0.9200 5.6550 1.0400 5.4150 1.0400 5.4150 0.6300 4.2550 0.6300
                 4.2550 0.4800 3.7750 0.4800 3.7750 0.9900 3.9350 0.9900 3.9350 1.1100 3.6550 1.1100
                 3.6550 0.3600 4.3750 0.3600 4.3750 0.5100 5.4150 0.5100 5.4150 0.3600 6.2350 0.3600
                 6.2350 0.7000 7.1850 0.7000 7.1850 1.3300 7.5150 1.3300 7.5150 0.4000 7.6350 0.4000 ;
        POLYGON  7.4950 2.2500 7.3750 2.2500 7.3750 2.0500 6.6650 2.0500 6.6650 2.2500 6.0150 2.2500
                 6.0150 2.0000 5.1350 2.0000 5.1350 2.2300 4.4950 2.2300 4.4950 1.5900 4.0150 1.5900
                 4.0150 2.2300 2.8850 2.2300 2.8850 1.6400 2.3250 1.6400 2.3250 2.2500 1.6750 2.2500
                 1.6750 1.5600 1.2350 1.5600 1.2350 1.6200 1.0950 1.6200 1.0950 1.7400 0.9750 1.7400
                 0.9750 1.4400 1.1150 1.4400 1.1150 1.0350 1.0950 1.0350 1.0950 0.6150 1.2150 0.6150
                 1.2150 0.9150 1.2350 0.9150 1.2350 1.4400 1.7950 1.4400 1.7950 2.1300 2.2050 2.1300
                 2.2050 1.5200 2.8850 1.5200 2.8850 1.0600 2.7950 1.0600 2.7950 0.9400 3.0350 0.9400
                 3.0350 1.0600 3.0050 1.0600 3.0050 2.1100 3.4150 2.1100 3.4150 1.1300 3.5350 1.1300
                 3.5350 2.1100 3.8950 2.1100 3.8950 1.4700 4.6150 1.4700 4.6150 2.1100 5.0150 2.1100
                 5.0150 1.8800 6.0150 1.8800 6.0150 1.1800 6.1350 1.1800 6.1350 2.1300 6.5450 2.1300
                 6.5450 1.9300 7.4950 1.9300 ;
        POLYGON  6.3750 2.0100 6.2550 2.0100 6.2550 1.0600 5.8950 1.0600 5.8950 1.2800 4.4150 1.2800
                 4.4150 1.3500 4.2950 1.3500 4.2950 1.1100 4.4150 1.1100 4.4150 1.1600 5.7750 1.1600
                 5.7750 0.7200 5.6550 0.7200 5.6550 0.6000 5.8950 0.6000 5.8950 0.9400 6.3750 0.9400 ;
        POLYGON  5.8950 1.7600 4.8950 1.7600 4.8950 1.9900 4.7750 1.9900 4.7750 1.6400 5.7750 1.6400
                 5.7750 1.5200 5.8950 1.5200 ;
        POLYGON  5.2950 1.0400 5.0550 1.0400 5.0550 0.9900 4.1750 0.9900 4.1750 1.3500 3.7750 1.3500
                 3.7750 1.9900 3.6550 1.9900 3.6550 1.2300 4.0550 1.2300 4.0550 0.8700 3.8950 0.8700
                 3.8950 0.6000 4.1350 0.6000 4.1350 0.7500 4.1750 0.7500 4.1750 0.8700 5.1750 0.8700
                 5.1750 0.9200 5.2950 0.9200 ;
        POLYGON  3.2950 1.9900 3.1750 1.9900 3.1750 0.8200 1.8550 0.8200 1.8550 1.0800 1.6550 1.0800
                 1.6550 0.8400 1.7350 0.8400 1.7350 0.7000 3.1750 0.7000 3.1750 0.5000 3.2950 0.5000 ;
        POLYGON  2.6750 1.0600 2.0950 1.0600 2.0950 1.4000 2.0350 1.4000 2.0350 2.0100 1.9150 2.0100
                 1.9150 1.3200 1.4150 1.3200 1.4150 0.4950 0.9750 0.4950 0.9750 1.0350 0.4750 1.0350
                 0.4750 1.2200 0.3550 1.2200 0.3550 0.9150 0.8550 0.9150 0.8550 0.3750 1.6150 0.3750
                 1.6150 0.7200 1.5350 0.7200 1.5350 1.2000 1.9750 1.2000 1.9750 0.9400 2.6750 0.9400 ;
    END
END DFFRHQX1

MACRO DFFQXL
    CLASS CORE ;
    FOREIGN DFFQXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6400 1.4650 0.8550 1.7250 ;
        RECT  0.6650 1.3850 0.8550 1.7250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9650 1.4900 5.2700 1.6650 ;
        RECT  4.8900 1.5200 5.2050 1.7200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9650 ;
        RECT  0.0700 1.4650 0.2550 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.0250 0.6700 5.2650 0.7900 ;
        RECT  5.0250 -0.1800 5.1450 0.7900 ;
        RECT  3.6050 0.4300 3.8450 0.5500 ;
        RECT  3.6050 -0.1800 3.7250 0.5500 ;
        RECT  1.9050 -0.1800 2.0250 0.8600 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1050 1.8700 5.2250 2.7900 ;
        RECT  3.5050 2.2900 3.7450 2.7900 ;
        RECT  1.7850 2.2900 2.0250 2.7900 ;
        RECT  0.5550 1.8450 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.6850 1.5100 5.6450 1.5100 5.6450 1.9900 5.5250 1.9900 5.5250 1.3900 5.5650 1.3900
                 5.5650 1.0300 4.7850 1.0300 4.7850 0.5000 4.0850 0.5000 4.0850 0.7900 3.3650 0.7900
                 3.3650 0.5000 3.0050 0.5000 3.0050 1.1500 3.2050 1.1500 3.2050 1.2700 2.6650 1.2700
                 2.6650 1.5300 2.5850 1.5300 2.5850 1.6500 2.4650 1.6500 2.4650 1.4100 2.5450 1.4100
                 2.5450 1.1500 2.8850 1.1500 2.8850 0.3800 3.4850 0.3800 3.4850 0.6700 3.9650 0.6700
                 3.9650 0.3800 4.1650 0.3800 4.1650 0.3600 4.4050 0.3600 4.4050 0.3800 4.9050 0.3800
                 4.9050 0.9100 5.5650 0.9100 5.5650 0.6200 5.6850 0.6200 ;
        POLYGON  5.4450 1.2700 5.3250 1.2700 5.3250 1.3700 4.7850 1.3700 4.7850 1.4000 4.6850 1.4000
                 4.6850 2.1700 2.9050 2.1700 2.9050 2.2500 2.1450 2.2500 2.1450 2.1700 0.9750 2.1700
                 0.9750 1.7250 1.0350 1.7250 1.0350 0.6800 1.1550 0.6800 1.1550 1.8450 1.0950 1.8450
                 1.0950 2.0500 2.2650 2.0500 2.2650 2.1300 2.7850 2.1300 2.7850 1.5500 2.8250 1.5500
                 2.8250 1.4300 2.9450 1.4300 2.9450 1.6700 2.9050 1.6700 2.9050 2.0500 4.5650 2.0500
                 4.5650 1.6500 4.1050 1.6500 4.1050 1.4100 4.2250 1.4100 4.2250 1.5300 4.5650 1.5300
                 4.5650 1.2500 4.6650 1.2500 4.6650 1.1600 4.7850 1.1600 4.7850 1.2500 5.2050 1.2500
                 5.2050 1.1500 5.4450 1.1500 ;
        POLYGON  4.5050 0.8600 4.3250 0.8600 4.3250 1.2900 3.9850 1.2900 3.9850 1.7700 4.3250 1.7700
                 4.3250 1.8100 4.4450 1.8100 4.4450 1.9300 4.2050 1.9300 4.2050 1.8900 3.8650 1.8900
                 3.8650 1.5000 3.6850 1.5000 3.6850 1.6200 3.5650 1.6200 3.5650 1.3800 3.8650 1.3800
                 3.8650 1.1700 4.2050 1.1700 4.2050 0.7400 4.3850 0.7400 4.3850 0.6200 4.5050 0.6200 ;
        POLYGON  3.7450 1.2600 3.4450 1.2600 3.4450 1.9300 3.0250 1.9300 3.0250 1.8100 3.3250 1.8100
                 3.3250 1.0300 3.1250 1.0300 3.1250 0.6200 3.2450 0.6200 3.2450 0.9100 3.4450 0.9100
                 3.4450 1.1400 3.6250 1.1400 3.6250 1.0200 3.7450 1.0200 ;
        POLYGON  2.7650 0.8000 2.3450 0.8000 2.3450 1.7700 2.6650 1.7700 2.6650 2.0100 2.5450 2.0100
                 2.5450 1.8900 2.2250 1.8900 2.2250 1.6500 1.7450 1.6500 1.7450 1.4100 1.8650 1.4100
                 1.8650 1.5300 2.2250 1.5300 2.2250 0.6800 2.7650 0.6800 ;
        POLYGON  2.1050 1.3100 1.9850 1.3100 1.9850 1.2900 1.6050 1.2900 1.6050 1.9300 1.3050 1.9300
                 1.3050 1.8100 1.4850 1.8100 1.4850 0.5600 0.9150 0.5600 0.9150 1.1600 0.5150 1.1600
                 0.5150 1.2800 0.3950 1.2800 0.3950 1.0400 0.7950 1.0400 0.7950 0.4400 1.6050 0.4400
                 1.6050 1.1700 1.9850 1.1700 1.9850 1.0700 2.1050 1.0700 ;
    END
END DFFQXL

MACRO DFFQX4
    CLASS CORE ;
    FOREIGN DFFQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9950 0.7200 2.2350 0.8400 ;
        RECT  2.0750 1.2800 2.1950 2.1100 ;
        RECT  2.0350 0.7200 2.1550 1.4000 ;
        RECT  1.2300 1.0250 2.1550 1.1450 ;
        RECT  1.2300 0.8850 1.3800 1.1450 ;
        RECT  1.2350 0.7200 1.3550 2.1100 ;
        RECT  1.2300 0.7200 1.3550 1.1450 ;
        RECT  1.0350 0.7200 1.3550 0.8400 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0600 0.5100 1.4350 ;
        RECT  0.3750 0.8400 0.4950 1.4350 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3950 1.2300 6.6550 1.4600 ;
        RECT  6.4550 1.1000 6.5750 1.5100 ;
        END
    END D
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.6750 -0.1800 6.7950 0.7400 ;
        RECT  5.0950 -0.1800 5.3350 0.3600 ;
        RECT  3.5550 -0.1800 3.6750 0.3800 ;
        RECT  2.4750 -0.1800 2.7150 0.3600 ;
        RECT  1.5150 -0.1800 1.7550 0.3600 ;
        RECT  0.5550 -0.1800 0.6750 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.5750 1.8700 6.6950 2.7900 ;
        RECT  4.9950 2.2900 5.2350 2.7900 ;
        RECT  3.3350 1.7500 3.4550 2.7900 ;
        RECT  2.4950 1.5900 2.6150 2.7900 ;
        RECT  1.6550 1.4600 1.7750 2.7900 ;
        RECT  0.8150 1.4600 0.9350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.3350 0.8400 7.2550 0.8400 7.2550 1.4200 7.1150 1.4200 7.1150 1.9900 6.9950 1.9900
                 6.9950 1.7500 6.1950 1.7500 6.1950 2.1700 4.2750 2.1700 4.2750 1.6500 3.9750 1.6500
                 3.9750 1.4100 4.0950 1.4100 4.0950 1.5300 4.5150 1.5300 4.5150 1.0000 4.6350 1.0000
                 4.6350 1.6500 4.3950 1.6500 4.3950 2.0500 6.0750 2.0500 6.0750 1.4300 6.1950 1.4300
                 6.1950 1.6300 6.9950 1.6300 6.9950 1.3000 7.1350 1.3000 7.1350 0.8400 7.0950 0.8400
                 7.0950 0.7200 7.3350 0.7200 ;
        POLYGON  7.0150 1.1800 6.7750 1.1800 6.7750 0.9800 6.2550 0.9800 6.2550 1.2400 6.1350 1.2400
                 6.1350 0.5400 5.7250 0.5400 5.7250 0.6000 5.7150 0.6000 5.7150 1.6500 5.5950 1.6500
                 5.5950 0.6000 4.8100 0.6000 4.8100 0.5400 4.1150 0.5400 4.1150 0.6200 3.3150 0.6200
                 3.3150 0.6000 0.9150 0.6000 0.9150 0.6600 0.2550 0.6600 0.2550 0.9000 0.2400 0.9000
                 0.2400 1.5550 0.5150 1.5550 0.5150 1.7950 0.3950 1.7950 0.3950 1.6750 0.1200 1.6750
                 0.1200 0.7800 0.1350 0.7800 0.1350 0.5400 0.7950 0.5400 0.7950 0.4800 3.4350 0.4800
                 3.4350 0.5000 3.9950 0.5000 3.9950 0.4000 4.2350 0.4000 4.2350 0.4200 4.9300 0.4200
                 4.9300 0.4800 5.6050 0.4800 5.6050 0.4200 6.2550 0.4200 6.2550 0.8600 6.8950 0.8600
                 6.8950 1.0600 7.0150 1.0600 ;
        POLYGON  6.0150 1.3100 5.9550 1.3100 5.9550 1.9300 5.7150 1.9300 5.7150 1.8900 5.3550 1.8900
                 5.3550 1.5900 4.9950 1.5900 4.9950 1.4700 5.4750 1.4700 5.4750 1.7700 5.8350 1.7700
                 5.8350 1.1900 5.8950 1.1900 5.8950 0.6600 6.0150 0.6600 ;
        POLYGON  5.3950 1.2900 4.8750 1.2900 4.8750 1.9300 4.5150 1.9300 4.5150 1.8100 4.7550 1.8100
                 4.7550 0.8400 4.6150 0.8400 4.6150 0.7200 4.8750 0.7200 4.8750 1.1700 5.2750 1.1700
                 5.2750 1.0500 5.3950 1.0500 ;
        POLYGON  4.3750 1.2900 3.8550 1.2900 3.8550 1.7700 4.0350 1.7700 4.0350 1.8100 4.1550 1.8100
                 4.1550 1.9300 3.9150 1.9300 3.9150 1.8900 3.7350 1.8900 3.7350 1.4900 3.1750 1.4900
                 3.1750 1.2500 3.2950 1.2500 3.2950 1.3700 3.7350 1.3700 3.7350 1.1700 4.2550 1.1700
                 4.2550 0.6600 4.3750 0.6600 ;
        POLYGON  3.6150 1.2500 3.4950 1.2500 3.4950 1.1300 3.0350 1.1300 3.0350 2.1100 2.9150 2.1100
                 2.9150 1.1300 2.5150 1.1300 2.5150 1.1600 2.2750 1.1600 2.2750 1.0100 3.0750 1.0100
                 3.0750 0.8400 2.9550 0.8400 2.9550 0.7200 3.1950 0.7200 3.1950 1.0100 3.6150 1.0100 ;
    END
END DFFQX4

MACRO DFFQX2
    CLASS CORE ;
    FOREIGN DFFQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1950 0.9250 0.4350 1.1650 ;
        RECT  0.0700 0.8850 0.3300 1.1450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4250 1.3150 1.5450 1.5550 ;
        RECT  1.2300 1.3150 1.5450 1.4350 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0650 0.6800 5.1850 1.6600 ;
        RECT  4.9650 1.5400 5.0850 2.1900 ;
        RECT  5.0000 1.1750 5.1850 1.6600 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.5450 -0.1800 5.6650 0.7600 ;
        RECT  4.5850 -0.1800 4.7050 0.7300 ;
        RECT  2.8450 -0.1800 2.9650 0.8900 ;
        RECT  1.4850 -0.1800 1.6050 0.3800 ;
        RECT  0.1350 -0.1800 0.2550 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.3850 1.5400 5.5050 2.7900 ;
        RECT  4.5450 1.8300 4.6650 2.7900 ;
        RECT  2.7850 2.1800 3.0250 2.3000 ;
        RECT  2.7850 2.1800 2.9050 2.7900 ;
        RECT  1.2650 1.9500 1.3850 2.7900 ;
        RECT  0.1350 1.4600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.1050 1.4200 5.9250 1.4200 5.9250 2.0600 5.8050 2.0600 5.8050 1.4200 5.3050 1.4200
                 5.3050 1.1800 5.4250 1.1800 5.4250 1.3000 5.9850 1.3000 5.9850 0.6200 6.1050 0.6200 ;
        POLYGON  5.8650 1.1800 5.7450 1.1800 5.7450 1.0000 5.3050 1.0000 5.3050 0.5600 4.9450 0.5600
                 4.9450 0.9700 3.9250 0.9700 3.9250 1.8900 4.0450 1.8900 4.0450 2.0100 3.8050 2.0100
                 3.8050 0.7200 4.0650 0.7200 4.0650 0.8500 4.8250 0.8500 4.8250 0.4400 5.4250 0.4400
                 5.4250 0.8800 5.8650 0.8800 ;
        POLYGON  4.2850 2.2500 3.1450 2.2500 3.1450 2.0600 2.6600 2.0600 2.6600 2.2500 1.7450 2.2500
                 1.7450 1.7950 1.1100 1.7950 1.1100 1.9150 0.9650 1.9150 0.9650 2.0900 0.8450 2.0900
                 0.8450 1.7950 0.9900 1.7950 0.9900 0.8400 0.8850 0.8400 0.8850 0.7200 1.1250 0.7200
                 1.1250 0.8400 1.1100 0.8400 1.1100 1.6750 1.7450 1.6750 1.7450 1.4900 1.8650 1.4900
                 1.8650 2.1300 2.5400 2.1300 2.5400 1.9400 3.2650 1.9400 3.2650 2.1300 4.1650 2.1300
                 4.1650 1.7500 4.0450 1.7500 4.0450 1.5100 4.1650 1.5100 4.1650 1.6300 4.2850 1.6300 ;
        POLYGON  4.2250 0.5000 3.7350 0.5000 3.7350 0.5400 3.6850 0.5400 3.6850 1.5800 3.5650 1.5800
                 3.5650 0.5400 3.2050 0.5400 3.2050 1.1300 2.4650 1.1300 2.4650 1.5800 2.2250 1.5800
                 2.2250 1.4600 2.3450 1.4600 2.3450 1.0100 2.4450 1.0100 2.4450 0.6000 1.8450 0.6000
                 1.8450 0.6200 1.2450 0.6200 1.2450 0.6000 0.6750 0.6000 0.6750 1.5800 0.5550 1.5800
                 0.5550 0.4800 1.0650 0.4800 1.0650 0.3800 1.3650 0.3800 1.3650 0.5000 1.7250 0.5000
                 1.7250 0.4800 1.9250 0.4800 1.9250 0.3800 2.1650 0.3800 2.1650 0.4800 2.5650 0.4800
                 2.5650 1.0100 3.0850 1.0100 3.0850 0.4200 3.6150 0.4200 3.6150 0.3800 4.2250 0.3800 ;
        POLYGON  3.6250 2.0100 3.3850 2.0100 3.3850 1.8200 3.3250 1.8200 3.3250 1.3700 2.5850 1.3700
                 2.5850 1.2500 3.3250 1.2500 3.3250 0.6600 3.4450 0.6600 3.4450 1.7000 3.5050 1.7000
                 3.5050 1.8900 3.6250 1.8900 ;
        POLYGON  3.1850 1.8200 2.3250 1.8200 2.3250 2.0100 1.9850 2.0100 1.9850 0.7200 2.3250 0.7200
                 2.3250 0.8400 2.1050 0.8400 2.1050 1.7000 3.0650 1.7000 3.0650 1.4900 3.1850 1.4900 ;
    END
END DFFQX2

MACRO DFFQX1
    CLASS CORE ;
    FOREIGN DFFQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.4550 0.9150 1.7250 ;
        RECT  0.6500 1.4400 0.8000 1.7250 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9850 1.4900 5.2250 1.7250 ;
        RECT  4.9450 1.4950 5.2050 1.7500 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 2.2050 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.1850 0.6800 5.4250 0.8000 ;
        RECT  5.1850 -0.1800 5.3050 0.8000 ;
        RECT  3.6250 0.4500 3.8650 0.5700 ;
        RECT  3.7450 -0.1800 3.8650 0.5700 ;
        RECT  1.9250 -0.1800 2.0450 0.8600 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1850 1.8700 5.3050 2.7900 ;
        RECT  3.5250 2.2900 3.7650 2.7900 ;
        RECT  1.8050 2.2900 2.0450 2.7900 ;
        RECT  0.5550 1.8450 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.8050 1.6100 5.7250 1.6100 5.7250 1.9900 5.6050 1.9900 5.6050 1.4900 5.6850 1.4900
                 5.6850 1.0400 4.8700 1.0400 4.8700 0.5000 4.1050 0.5000 4.1050 0.8100 3.3850 0.8100
                 3.3850 0.5000 3.0250 0.5000 3.0250 1.1700 3.2250 1.1700 3.2250 1.2900 2.6650 1.2900
                 2.6650 1.5300 2.5850 1.5300 2.5850 1.6500 2.4650 1.6500 2.4650 1.4100 2.5450 1.4100
                 2.5450 1.1700 2.9050 1.1700 2.9050 0.3800 3.5050 0.3800 3.5050 0.6900 3.9850 0.6900
                 3.9850 0.3800 4.2650 0.3800 4.2650 0.3600 4.5050 0.3600 4.5050 0.3800 4.9900 0.3800
                 4.9900 0.9200 5.6650 0.9200 5.6650 0.6200 5.7850 0.6200 5.7850 0.7400 5.8050 0.7400 ;
        POLYGON  5.5650 1.3700 4.8050 1.3700 4.8050 1.4100 4.7050 1.4100 4.7050 2.1700 2.9250 2.1700
                 2.9250 2.2500 2.2750 2.2500 2.2750 2.1700 0.9750 2.1700 0.9750 1.8450 1.0350 1.8450
                 1.0350 0.6800 1.1550 0.6800 1.1550 2.0500 2.3950 2.0500 2.3950 2.1300 2.8050 2.1300
                 2.8050 1.6100 2.7850 1.6100 2.7850 1.4900 3.0250 1.4900 3.0250 1.6100 2.9250 1.6100
                 2.9250 2.0500 4.5850 2.0500 4.5850 1.6500 4.1250 1.6500 4.1250 1.4100 4.2450 1.4100
                 4.2450 1.5300 4.5850 1.5300 4.5850 1.2500 4.6850 1.2500 4.6850 1.1700 4.8050 1.1700
                 4.8050 1.2500 5.5650 1.2500 ;
        POLYGON  4.7250 1.0500 4.0050 1.0500 4.0050 1.7700 4.3450 1.7700 4.3450 1.8100 4.4650 1.8100
                 4.4650 1.9300 4.2250 1.9300 4.2250 1.8900 3.8850 1.8900 3.8850 1.4500 3.7050 1.4500
                 3.7050 1.5700 3.5850 1.5700 3.5850 1.3300 3.8850 1.3300 3.8850 0.9300 4.6050 0.9300
                 4.6050 0.6200 4.7250 0.6200 ;
        POLYGON  3.7650 1.2100 3.4650 1.2100 3.4650 1.9300 3.0450 1.9300 3.0450 1.8100 3.3450 1.8100
                 3.3450 1.0500 3.1450 1.0500 3.1450 0.6200 3.2650 0.6200 3.2650 0.9300 3.4650 0.9300
                 3.4650 1.0900 3.6450 1.0900 3.6450 0.9700 3.7650 0.9700 ;
        POLYGON  2.7850 0.8000 2.3450 0.8000 2.3450 1.7700 2.6850 1.7700 2.6850 2.0100 2.5650 2.0100
                 2.5650 1.8900 2.2250 1.8900 2.2250 1.5300 1.6450 1.5300 1.6450 1.4100 2.2250 1.4100
                 2.2250 0.6800 2.7850 0.6800 ;
        POLYGON  2.1050 1.2000 1.5250 1.2000 1.5250 1.8100 1.5650 1.8100 1.5650 1.9300 1.3250 1.9300
                 1.3250 1.8100 1.4050 1.8100 1.4050 0.7400 1.4250 0.7400 1.4250 0.5600 0.9150 0.5600
                 0.9150 0.9700 0.5350 0.9700 0.5350 1.2400 0.4150 1.2400 0.4150 0.8500 0.7950 0.8500
                 0.7950 0.4400 1.5450 0.4400 1.5450 0.8600 1.5250 0.8600 1.5250 1.0800 2.1050 1.0800 ;
    END
END DFFQX1

MACRO DFFNSRXL
    CLASS CORE ;
    FOREIGN DFFNSRXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9450 1.4850 2.0650 1.7500 ;
        RECT  1.8100 1.4450 1.9600 1.7250 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7550 2.1300 7.6350 2.2500 ;
        RECT  6.7550 1.7300 6.8750 2.2500 ;
        RECT  6.1550 1.7300 6.8750 1.8500 ;
        RECT  5.1850 1.8400 6.2750 1.9000 ;
        RECT  5.6950 1.7800 6.8750 1.8500 ;
        RECT  5.1850 1.8400 5.8150 1.9600 ;
        RECT  3.9150 1.7400 5.3050 1.8600 ;
        RECT  3.2150 1.8100 4.0350 1.9300 ;
        RECT  3.2150 1.2500 3.4550 1.3700 ;
        RECT  3.2150 1.2500 3.3350 1.9300 ;
        RECT  2.9150 1.5200 3.3350 1.6700 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3750 0.8700 9.5150 1.2200 ;
        RECT  9.3300 0.8100 9.5000 1.1600 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.4550 1.2000 10.7150 1.4300 ;
        RECT  10.4650 1.2000 10.5850 1.6100 ;
        END
    END CKN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.5800 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3650 1.5850 1.4850 2.0900 ;
        RECT  1.3650 0.6800 1.4850 0.9600 ;
        RECT  1.2300 1.4650 1.4450 1.7250 ;
        RECT  1.3250 0.8400 1.4450 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  10.7650 -0.1800 10.8850 0.4000 ;
        RECT  9.3550 -0.1800 9.4750 0.3800 ;
        RECT  8.0350 -0.1800 8.2750 0.3300 ;
        RECT  3.0750 -0.1800 3.3150 0.3200 ;
        RECT  1.7850 -0.1800 1.9050 0.9200 ;
        RECT  0.6150 -0.1800 0.7350 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  10.7050 1.6700 10.8250 2.7900 ;
        RECT  9.3150 1.9000 9.4350 2.7900 ;
        RECT  7.7750 2.1300 7.8950 2.7900 ;
        RECT  6.1750 2.2900 6.4150 2.7900 ;
        RECT  4.4150 2.2200 4.6550 2.7900 ;
        RECT  3.0750 2.2900 3.3150 2.7900 ;
        RECT  1.7850 1.9700 1.9050 2.7900 ;
        RECT  0.5550 1.4600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.4650 1.8500 10.2150 1.8500 10.2150 0.9600 10.2850 0.9600 10.2850 0.6000
                 9.7150 0.6000 9.7150 0.6200 9.1050 0.6200 9.1050 0.5700 7.5950 0.5700 7.5950 0.4800
                 7.4750 0.4800 7.4750 0.3600 7.7150 0.3600 7.7150 0.4500 8.5750 0.4500 8.5750 0.3800
                 8.8150 0.3800 8.8150 0.4500 9.2250 0.4500 9.2250 0.5000 9.5950 0.5000 9.5950 0.3800
                 9.9150 0.3800 9.9150 0.4800 10.4050 0.4800 10.4050 1.0800 10.3350 1.0800
                 10.3350 1.7300 10.4650 1.7300 ;
        POLYGON  10.0750 0.8400 9.9550 0.8400 9.9550 1.7800 9.8750 1.7800 9.8750 2.0200 9.7550 2.0200
                 9.7550 1.7800 9.0950 1.7800 9.0950 2.2000 8.3750 2.2000 8.3750 2.0100 6.9950 2.0100
                 6.9950 1.6100 6.6750 1.6100 6.6750 1.3500 6.2450 1.3500 6.2450 1.2300 6.7950 1.2300
                 6.7950 1.4900 7.1150 1.4900 7.1150 1.8900 8.4950 1.8900 8.4950 2.0800 8.9750 2.0800
                 8.9750 1.5300 8.5150 1.5300 8.5150 1.2900 8.6350 1.2900 8.6350 1.4100 8.9750 1.4100
                 8.9750 1.2800 9.2350 1.2800 9.2350 1.4000 9.0950 1.4000 9.0950 1.6600 9.8350 1.6600
                 9.8350 0.7200 10.0750 0.7200 ;
        POLYGON  8.9750 0.8400 8.8550 0.8400 8.8550 1.1300 8.3950 1.1300 8.3950 1.6500 8.7350 1.6500
                 8.7350 1.8400 8.8550 1.8400 8.8550 1.9600 8.6150 1.9600 8.6150 1.7700 8.2750 1.7700
                 8.2750 1.1300 7.1550 1.1300 7.1550 1.0100 8.7350 1.0100 8.7350 0.7200 8.9750 0.7200 ;
        POLYGON  8.1550 1.5300 7.9150 1.5300 7.9150 1.3700 7.3550 1.3700 7.3550 1.6500 7.4750 1.6500
                 7.4750 1.7700 7.2350 1.7700 7.2350 1.3700 6.9150 1.3700 6.9150 1.1100 6.1250 1.1100
                 6.1250 1.5800 6.0350 1.5800 6.0350 1.6600 5.7850 1.6600 5.7850 1.5400 5.9150 1.5400
                 5.9150 1.4600 6.0050 1.4600 6.0050 0.8600 5.8850 0.8600 5.8850 0.6200 6.0050 0.6200
                 6.0050 0.7400 6.1250 0.7400 6.1250 0.9900 6.9150 0.9900 6.9150 0.7500 6.9950 0.7500
                 6.9950 0.6300 7.1150 0.6300 7.1150 0.8700 7.0350 0.8700 7.0350 1.2500 8.0350 1.2500
                 8.0350 1.4100 8.1550 1.4100 ;
        POLYGON  7.5950 0.8100 7.3550 0.8100 7.3550 0.7200 7.2350 0.7200 7.2350 0.5100 6.6950 0.5100
                 6.6950 0.8700 6.5750 0.8700 6.5750 0.3900 7.3550 0.3900 7.3550 0.6000 7.4750 0.6000
                 7.4750 0.6900 7.5950 0.6900 ;
        POLYGON  6.6350 2.0900 6.5150 2.0900 6.5150 2.1400 6.0550 2.1400 6.0550 2.2000 4.8750 2.2000
                 4.8750 2.1000 4.2750 2.1000 4.2750 2.2200 4.1550 2.2200 4.1550 2.1700 2.2050 2.1700
                 2.2050 1.8500 2.2650 1.8500 2.2650 0.6800 2.3850 0.6800 2.3850 2.0500 4.1550 2.0500
                 4.1550 1.9800 4.9950 1.9800 4.9950 2.0800 5.9350 2.0800 5.9350 2.0200 6.3950 2.0200
                 6.3950 1.9700 6.6350 1.9700 ;
        POLYGON  5.8850 1.3400 5.6450 1.3400 5.6450 0.4800 5.2050 0.4800 5.2050 0.3600 5.7650 0.3600
                 5.7650 1.2200 5.8850 1.2200 ;
        POLYGON  5.5450 1.7200 5.4250 1.7200 5.4250 1.5800 5.4050 1.5800 5.4050 1.3800 3.5750 1.3800
                 3.5750 1.1300 3.0950 1.1300 3.0950 1.1800 2.8550 1.1800 2.8550 1.0600 2.9750 1.0600
                 2.9750 1.0100 3.6950 1.0100 3.6950 1.2600 5.4050 1.2600 5.4050 0.6200 5.5250 0.6200
                 5.5250 1.4600 5.5450 1.4600 ;
        POLYGON  5.1850 1.6200 3.7950 1.6200 3.7950 1.6900 3.5550 1.6900 3.5550 1.5700 3.6750 1.5700
                 3.6750 1.5000 5.1850 1.5000 ;
        POLYGON  5.1050 0.8600 4.9550 0.8600 4.9550 1.1400 4.3550 1.1400 4.3550 0.9000 4.1750 0.9000
                 4.1750 0.6600 4.2950 0.6600 4.2950 0.7800 4.4750 0.7800 4.4750 1.0200 4.8350 1.0200
                 4.8350 0.7400 4.9850 0.7400 4.9850 0.6200 5.1050 0.6200 ;
        POLYGON  4.7150 0.9000 4.5950 0.9000 4.5950 0.5400 4.0550 0.5400 4.0550 0.7600 3.7950 0.7600
                 3.7950 0.8400 3.5550 0.8400 3.5550 0.7200 3.6750 0.7200 3.6750 0.6400 3.9350 0.6400
                 3.9350 0.4200 4.7150 0.4200 ;
        POLYGON  3.8150 0.5200 3.5550 0.5200 3.5550 0.5600 2.7750 0.5600 2.7750 0.9000 2.7350 0.9000
                 2.7350 1.3000 2.7750 1.3000 2.7750 1.7500 2.6550 1.7500 2.6550 1.4200 2.6150 1.4200
                 2.6150 0.7800 2.6550 0.7800 2.6550 0.5600 2.1450 0.5600 2.1450 1.2000 1.5650 1.2000
                 1.5650 1.0800 2.0250 1.0800 2.0250 0.4400 3.4350 0.4400 3.4350 0.4000 3.8150 0.4000 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFNSRXL

MACRO DFFNSRX4
    CLASS CORE ;
    FOREIGN DFFNSRX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 13.6300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.3250 0.5100 1.7250 ;
        RECT  0.3900 1.2200 0.5100 1.7250 ;
        END
    END CKN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6300 1.4650 0.8400 1.7250 ;
        RECT  0.6550 1.3800 0.8400 1.7250 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 0.9450 4.2450 1.1450 ;
        RECT  3.7850 0.9200 4.0450 1.1450 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.5050 1.0900 5.0250 1.2100 ;
        RECT  4.3650 1.2300 4.6250 1.3800 ;
        RECT  4.5050 1.0900 4.6250 1.3800 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.4750 0.7400 10.6750 0.8600 ;
        RECT  10.3750 1.4200 10.4950 2.1900 ;
        RECT  10.1950 1.4200 10.4950 1.5400 ;
        RECT  9.5850 1.3000 10.3150 1.4200 ;
        RECT  9.5850 1.2300 9.8450 1.4200 ;
        RECT  9.5350 1.4200 9.8350 1.5400 ;
        RECT  9.7150 0.7400 9.8350 1.5400 ;
        RECT  9.5350 1.4200 9.6550 2.1900 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.3950 0.7400 12.5950 0.8600 ;
        RECT  12.0550 1.4200 12.1750 2.1900 ;
        RECT  11.8750 1.4200 12.1750 1.5400 ;
        RECT  11.0900 1.3000 11.9950 1.4200 ;
        RECT  11.2150 1.3000 11.5150 1.5400 ;
        RECT  11.3950 0.7400 11.5150 1.5400 ;
        RECT  11.2150 1.3000 11.3350 2.1900 ;
        RECT  11.0900 1.1750 11.2400 1.4350 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 13.6300 0.1800 ;
        RECT  12.9550 -0.1800 13.0750 0.7300 ;
        RECT  11.8750 -0.1800 12.1150 0.3800 ;
        RECT  10.9150 -0.1800 11.1550 0.3800 ;
        RECT  9.9550 -0.1800 10.1950 0.3800 ;
        RECT  8.9950 -0.1800 9.1150 0.8200 ;
        RECT  8.1550 -0.1800 8.2750 0.8600 ;
        RECT  4.6450 0.6100 4.8850 0.7300 ;
        RECT  4.7650 -0.1800 4.8850 0.7300 ;
        RECT  2.0950 -0.1800 2.3350 0.3200 ;
        RECT  0.5550 -0.1800 0.6750 0.8600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 13.6300 2.7900 ;
        RECT  12.4750 1.5400 12.5950 2.7900 ;
        RECT  11.6350 1.5400 11.7550 2.7900 ;
        RECT  10.7950 1.5400 10.9150 2.7900 ;
        RECT  9.9550 1.5400 10.0750 2.7900 ;
        RECT  9.1150 1.6400 9.2350 2.7900 ;
        RECT  8.2750 1.7000 8.3950 2.7900 ;
        RECT  7.1550 1.8800 7.3950 2.0000 ;
        RECT  7.1550 1.8800 7.2750 2.7900 ;
        RECT  3.9850 2.2200 4.2250 2.7900 ;
        RECT  2.8050 2.2250 3.0450 2.7900 ;
        RECT  1.8950 2.2250 2.0150 2.7900 ;
        RECT  0.5550 1.9200 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  13.4950 0.9200 13.3350 0.9200 13.3350 1.4200 13.0150 1.4200 13.0150 2.1900
                 12.8950 2.1900 12.8950 1.4200 12.2950 1.4200 12.2950 1.2800 12.5350 1.2800
                 12.5350 1.3000 13.2150 1.3000 13.2150 0.8000 13.3750 0.8000 13.3750 0.6800
                 13.4950 0.6800 ;
        POLYGON  13.0950 1.1800 12.8550 1.1800 12.8550 0.9700 12.7150 0.9700 12.7150 0.6200
                 9.3550 0.6200 9.3550 1.0600 8.8550 1.0600 8.8550 1.1800 9.4550 1.1800 9.4550 1.3000
                 8.8550 1.3000 8.8550 1.7600 8.8150 1.7600 8.8150 2.1600 8.6950 2.1600 8.6950 1.6400
                 8.7350 1.6400 8.7350 1.2200 7.6150 1.2200 7.6150 1.1000 8.5750 1.1000 8.5750 0.6800
                 8.6950 0.6800 8.6950 0.9400 9.2350 0.9400 9.2350 0.5000 12.8350 0.5000 12.8350 0.8500
                 12.9750 0.8500 12.9750 1.0600 13.0950 1.0600 ;
        POLYGON  8.6150 1.5200 6.2650 1.5200 6.2650 1.7100 6.0250 1.7100 6.0250 0.6700 6.1450 0.6700
                 6.1450 1.4000 8.3750 1.4000 8.3750 1.3600 8.6150 1.3600 ;
        POLYGON  8.0350 1.8800 7.5150 1.8800 7.5150 1.7600 6.4450 1.7600 6.4450 1.6400 7.6350 1.6400
                 7.6350 1.7600 8.0350 1.7600 ;
        POLYGON  7.8550 0.8600 7.7350 0.8600 7.7350 0.5600 7.0750 0.5600 7.0750 0.8000 6.8350 0.8000
                 6.8350 0.6800 6.9550 0.6800 6.9550 0.4400 7.8550 0.4400 ;
        POLYGON  7.4950 0.8000 7.3150 0.8000 7.3150 1.0400 6.5950 1.0400 6.5950 0.9100 6.5050 0.9100
                 6.5050 0.6700 6.6250 0.6700 6.6250 0.7900 6.7150 0.7900 6.7150 0.9200 7.1950 0.9200
                 7.1950 0.6800 7.4950 0.6800 ;
        POLYGON  7.2350 1.2800 6.3550 1.2800 6.3550 1.1500 6.2650 1.1500 6.2650 0.5500 5.3050 0.5500
                 5.3050 1.5300 5.0650 1.5300 5.0650 1.4100 5.1850 1.4100 5.1850 0.9700 4.3900 0.9700
                 4.3900 0.4800 4.0850 0.4800 4.0850 0.3600 4.5100 0.3600 4.5100 0.8500 5.1850 0.8500
                 5.1850 0.4300 6.3850 0.4300 6.3850 1.0300 6.4750 1.0300 6.4750 1.1600 7.2350 1.1600 ;
        POLYGON  7.0250 2.0500 6.7850 2.0500 6.7850 2.0100 4.5850 2.0100 4.5850 1.8600 3.7650 1.8600
                 3.7650 1.6250 2.7650 1.6250 2.7650 1.2200 2.8850 1.2200 2.8850 1.5050 3.8850 1.5050
                 3.8850 1.7400 4.7050 1.7400 4.7050 1.8900 5.7850 1.8900 5.7850 1.1700 5.6650 1.1700
                 5.6650 1.0500 5.9050 1.0500 5.9050 1.8900 6.9050 1.8900 6.9050 1.9300 7.0250 1.9300 ;
        POLYGON  6.0050 2.2500 4.3450 2.2500 4.3450 2.1000 3.5250 2.1000 3.5250 1.8650 2.4350 1.8650
                 2.4350 1.7450 2.5250 1.7450 2.5250 1.4600 1.5350 1.4600 1.5350 1.3200 1.7750 1.3200
                 1.7750 1.3400 2.5250 1.3400 2.5250 0.7200 2.7650 0.7200 2.7650 0.8400 2.6450 0.8400
                 2.6450 1.7450 3.6450 1.7450 3.6450 1.9800 4.4650 1.9800 4.4650 2.1300 6.0050 2.1300 ;
        POLYGON  5.7250 0.9300 5.5450 0.9300 5.5450 1.5300 5.6650 1.5300 5.6650 1.7700 4.8250 1.7700
                 4.8250 1.6200 4.0050 1.6200 4.0050 1.3850 3.5450 1.3850 3.5450 1.1000 2.8850 1.1000
                 2.8850 0.5600 1.8550 0.5600 1.8550 0.4800 1.7350 0.4800 1.7350 0.3600 1.9750 0.3600
                 1.9750 0.4400 3.0050 0.4400 3.0050 0.9800 3.5450 0.9800 3.5450 0.8000 3.4850 0.8000
                 3.4850 0.6800 3.7250 0.6800 3.7250 0.8000 3.6650 0.8000 3.6650 1.2650 4.2450 1.2650
                 4.2450 1.5000 4.9450 1.5000 4.9450 1.6500 5.4250 1.6500 5.4250 0.8100 5.6050 0.8100
                 5.6050 0.6700 5.7250 0.6700 ;
        POLYGON  4.1650 0.8000 3.8450 0.8000 3.8450 0.5600 3.3650 0.5600 3.3650 0.6200 3.2450 0.6200
                 3.2450 0.8600 3.1250 0.8600 3.1250 0.5000 3.2450 0.5000 3.2450 0.4400 3.9650 0.4400
                 3.9650 0.6800 4.1650 0.6800 ;
        POLYGON  3.4050 2.2500 3.1650 2.2500 3.1650 2.1050 1.1950 2.1050 1.1950 1.8400 1.2950 1.8400
                 1.2950 0.9600 1.2550 0.9600 1.2550 0.6200 1.3750 0.6200 1.3750 0.8400 1.4150 0.8400
                 1.4150 1.9850 3.2850 1.9850 3.2850 2.1300 3.4050 2.1300 ;
        POLYGON  2.4050 1.2200 2.2850 1.2200 2.2850 1.0600 1.6950 1.0600 1.6950 1.1800 1.5750 1.1800
                 1.5750 0.7200 1.4950 0.7200 1.4950 0.5000 1.1350 0.5000 1.1350 1.4800 1.1750 1.4800
                 1.1750 1.7200 1.0150 1.7200 1.0150 1.1000 0.2400 1.1000 0.2400 1.8450 0.2550 1.8450
                 0.2550 2.0850 0.1350 2.0850 0.1350 1.9650 0.1200 1.9650 0.1200 0.8600 0.1350 0.8600
                 0.1350 0.6200 0.2550 0.6200 0.2550 0.9800 1.0150 0.9800 1.0150 0.3800 1.6150 0.3800
                 1.6150 0.6000 1.6950 0.6000 1.6950 0.9400 2.4050 0.9400 ;
    END
END DFFNSRX4

MACRO DFFNSRX2
    CLASS CORE ;
    FOREIGN DFFNSRX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.6000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4100 1.3450 0.5300 1.8000 ;
        RECT  0.3600 1.2900 0.5100 1.7250 ;
        END
    END CKN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3650 1.1650 4.6250 1.3800 ;
        RECT  4.4650 1.0000 4.5850 1.3800 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0000 1.0300 5.1500 1.4350 ;
        RECT  4.9850 1.0000 5.1050 1.4100 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.4600 0.8700 1.7800 ;
        RECT  0.6500 1.4550 0.8000 1.7800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.5650 1.4650 9.7900 1.7250 ;
        RECT  9.5650 1.3400 9.7600 1.7250 ;
        RECT  9.6200 0.5900 9.7400 1.7250 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5100 1.4650 10.6600 1.7250 ;
        RECT  10.4800 1.4500 10.6450 1.5700 ;
        RECT  10.4800 0.7100 10.6000 1.5700 ;
        RECT  10.4600 0.5900 10.5800 0.8300 ;
        END
    END QN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.6000 0.1800 ;
        RECT  10.8800 -0.1800 11.0000 0.6400 ;
        RECT  10.0400 -0.1800 10.1600 0.6400 ;
        RECT  9.2000 -0.1800 9.3200 0.7300 ;
        RECT  7.0700 -0.1800 7.1900 0.7800 ;
        RECT  4.6050 0.4800 4.8450 0.6400 ;
        RECT  4.6050 -0.1800 4.7250 0.6400 ;
        RECT  2.1500 -0.1800 2.3900 0.3200 ;
        RECT  0.6700 -0.1800 0.7900 0.8600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.6000 2.7900 ;
        RECT  11.0050 2.0850 11.1250 2.7900 ;
        RECT  10.0450 2.0850 10.1650 2.7900 ;
        RECT  9.0850 1.8600 9.2050 2.7900 ;
        RECT  7.9700 1.8700 8.3100 1.9900 ;
        RECT  8.1900 1.6300 8.3100 1.9900 ;
        RECT  7.9700 1.8700 8.0900 2.7900 ;
        RECT  7.1300 1.8600 7.2500 2.7900 ;
        RECT  4.1900 2.2750 4.4300 2.7900 ;
        RECT  3.0050 2.1000 3.1250 2.7900 ;
        RECT  2.1900 2.1000 2.3100 2.7900 ;
        RECT  0.5900 1.9200 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  11.4650 1.5800 11.3450 1.5800 11.3450 0.8800 10.8400 0.8800 10.8400 1.1700
                 10.7200 1.1700 10.7200 0.7600 11.3000 0.7600 11.3000 0.4000 11.4200 0.4000
                 11.4200 0.7600 11.4650 0.7600 ;
        POLYGON  11.1600 1.9650 9.3250 1.9650 9.3250 1.7400 8.7250 1.7400 8.7250 2.2500 8.2100 2.2500
                 8.2100 2.1300 8.6050 2.1300 8.6050 1.6200 9.3050 1.6200 9.3050 1.0100 8.7800 1.0100
                 8.7800 0.5900 8.9000 0.5900 8.9000 0.8900 9.4250 0.8900 9.4250 1.6200 9.4450 1.6200
                 9.4450 1.8450 9.9100 1.8450 9.9100 1.2600 9.9000 1.2600 9.9000 1.0200 10.0300 1.0200
                 10.0300 1.8450 11.0400 1.8450 11.0400 1.0000 11.1600 1.0000 ;
        POLYGON  8.8850 1.5000 6.3200 1.5000 6.3200 1.7700 6.2000 1.7700 6.2000 0.6700 6.3200 0.6700
                 6.3200 1.3800 8.7650 1.3800 8.7650 1.1300 8.8850 1.1300 ;
        POLYGON  8.5100 1.0200 7.6000 1.0200 7.6000 0.8400 7.5500 0.8400 7.5500 0.6000 7.6700 0.6000
                 7.6700 0.7200 7.7200 0.7200 7.7200 0.9000 8.3900 0.9000 8.3900 0.6000 8.5100 0.6000 ;
        POLYGON  8.2300 1.2600 6.4400 1.2600 6.4400 0.5500 5.2650 0.5500 5.2650 0.7600 5.3900 0.7600
                 5.3900 1.4100 5.5100 1.4100 5.5100 1.5300 5.2700 1.5300 5.2700 0.8800 4.3050 0.8800
                 4.3050 0.4800 4.0650 0.4800 4.0650 0.3600 4.4250 0.3600 4.4250 0.7600 4.9650 0.7600
                 4.9650 0.6400 5.1450 0.6400 5.1450 0.4300 6.5600 0.4300 6.5600 1.1400 8.2300 1.1400 ;
        POLYGON  8.1500 0.7800 7.9100 0.7800 7.9100 0.6600 7.8400 0.6600 7.8400 0.4800 7.4300 0.4800
                 7.4300 1.0200 6.6800 1.0200 6.6800 0.6700 6.8000 0.6700 6.8000 0.9000 7.3100 0.9000
                 7.3100 0.3600 7.9600 0.3600 7.9600 0.5400 8.0300 0.5400 8.0300 0.6600 8.1500 0.6600 ;
        POLYGON  7.6700 1.9800 7.5500 1.9800 7.5500 1.8600 7.3700 1.8600 7.3700 1.7400 6.5600 1.7400
                 6.5600 1.6200 7.4900 1.6200 7.4900 1.7400 7.6700 1.7400 ;
        POLYGON  6.5200 2.1500 6.2200 2.1500 6.2200 2.0100 4.7900 2.0100 4.7900 1.9150 3.8850 1.9150
                 3.8850 1.3600 2.8100 1.3600 2.8100 1.2400 4.0050 1.2400 4.0050 1.7950 4.9100 1.7950
                 4.9100 1.8900 5.9600 1.8900 5.9600 1.2300 5.9000 1.2300 5.9000 0.9900 6.0200 0.9900
                 6.0200 1.1100 6.0800 1.1100 6.0800 1.8900 6.3400 1.8900 6.3400 2.0300 6.5200 2.0300 ;
        POLYGON  6.1000 2.2500 4.5500 2.2500 4.5500 2.1550 3.6450 2.1550 3.6450 2.0100 3.4850 2.0100
                 3.4850 1.7400 2.5500 1.7400 2.5500 1.4400 1.5700 1.4400 1.5700 1.3200 2.5700 1.3200
                 2.5700 0.9200 2.5500 0.9200 2.5500 0.6800 2.6700 0.6800 2.6700 0.8000 2.6900 0.8000
                 2.6900 1.6200 3.6050 1.6200 3.6050 1.8900 3.7650 1.8900 3.7650 2.0350 4.6700 2.0350
                 4.6700 2.1300 6.1000 2.1300 ;
        POLYGON  5.8400 1.7700 5.0300 1.7700 5.0300 1.6750 4.1250 1.6750 4.1250 1.1200 2.9250 1.1200
                 2.9250 0.5600 1.9100 0.5600 1.9100 0.4800 1.7900 0.4800 1.7900 0.3600 2.0300 0.3600
                 2.0300 0.4400 3.0450 0.4400 3.0450 1.0000 3.5850 1.0000 3.5850 0.6400 3.7050 0.6400
                 3.7050 1.0000 4.2450 1.0000 4.2450 1.5000 4.3650 1.5000 4.3650 1.5550 5.1500 1.5550
                 5.1500 1.6500 5.6600 1.6500 5.6600 0.6700 5.7800 0.6700 5.7800 1.5300 5.8400 1.5300 ;
        POLYGON  4.1850 0.8200 3.8250 0.8200 3.8250 0.5200 3.4650 0.5200 3.4650 0.6400 3.2850 0.6400
                 3.2850 0.8800 3.1650 0.8800 3.1650 0.5200 3.3450 0.5200 3.3450 0.4000 3.9450 0.4000
                 3.9450 0.7000 4.1850 0.7000 ;
        POLYGON  3.5250 2.2500 3.2450 2.2500 3.2450 1.9800 1.4500 1.9800 1.4500 2.0400 1.3300 2.0400
                 1.3300 1.3600 1.3100 1.3600 1.3100 0.6200 1.4300 0.6200 1.4300 1.2400 1.4500 1.2400
                 1.4500 1.8600 3.3650 1.8600 3.3650 2.1300 3.5250 2.1300 ;
        POLYGON  2.4500 1.1800 1.5700 1.1800 1.5700 0.9400 1.5500 0.9400 1.5500 0.5000 1.1900 0.5000
                 1.1900 1.4800 1.2100 1.4800 1.2100 1.7200 1.0700 1.7200 1.0700 1.1700 0.2400 1.1700
                 0.2400 1.8450 0.2900 1.8450 0.2900 2.0850 0.1700 2.0850 0.1700 1.9650 0.1200 1.9650
                 0.1200 0.7400 0.2500 0.7400 0.2500 0.6200 0.3700 0.6200 0.3700 0.8600 0.2400 0.8600
                 0.2400 1.0500 1.0700 1.0500 1.0700 0.3800 1.6700 0.3800 1.6700 0.8200 1.6900 0.8200
                 1.6900 1.0000 1.8100 1.0000 1.8100 1.0600 2.4500 1.0600 ;
    END
END DFFNSRX2

MACRO DFFNSRX1
    CLASS CORE ;
    FOREIGN DFFNSRX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.3100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9050 1.2100 2.1450 1.4400 ;
        RECT  1.7550 1.2300 2.0150 1.4850 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7950 2.1300 7.6750 2.2500 ;
        RECT  6.7950 1.7800 6.9150 2.2500 ;
        RECT  5.5950 1.7800 6.9150 1.9000 ;
        RECT  5.1150 1.8400 5.7150 1.9600 ;
        RECT  5.1150 1.7000 5.2350 1.9600 ;
        RECT  4.0050 1.7000 5.2350 1.8200 ;
        RECT  3.2550 1.7700 4.1250 1.8900 ;
        RECT  3.2550 1.5200 3.4650 1.8900 ;
        RECT  3.2550 1.0000 3.3750 1.8900 ;
        RECT  3.2050 1.5200 3.4650 1.6700 ;
        RECT  3.1350 1.0000 3.3750 1.1200 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.4350 0.8350 9.7900 1.2100 ;
        RECT  9.4350 0.8350 9.5550 1.2200 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.5100 0.8650 10.6600 1.3200 ;
        RECT  10.5200 0.8650 10.6400 1.3400 ;
        END
    END CKN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.6800 0.2550 1.9900 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3850 1.4900 1.5050 2.1400 ;
        RECT  1.3650 0.6100 1.4850 0.8500 ;
        RECT  1.2300 1.4650 1.4250 1.7250 ;
        RECT  1.3050 0.7300 1.4250 1.7250 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.3100 0.1800 ;
        RECT  10.7800 -0.1800 10.9000 0.7450 ;
        RECT  9.4300 -0.1800 9.5500 0.3800 ;
        RECT  8.0750 -0.1800 8.3150 0.3600 ;
        RECT  3.0750 -0.1800 3.3150 0.3200 ;
        RECT  1.7850 -0.1800 1.9050 0.8500 ;
        RECT  0.5550 -0.1800 0.6750 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.3100 2.7900 ;
        RECT  10.7800 1.4600 10.9000 2.7900 ;
        RECT  9.3550 1.9000 9.4750 2.7900 ;
        RECT  7.8150 2.1300 7.9350 2.7900 ;
        RECT  6.0750 2.2600 6.3150 2.7900 ;
        RECT  4.4850 2.1800 4.7250 2.3000 ;
        RECT  4.4850 2.1800 4.6050 2.7900 ;
        RECT  3.1650 2.2500 3.4050 2.7900 ;
        RECT  1.8050 1.6050 1.9250 2.7900 ;
        RECT  0.5550 1.3400 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.4800 0.7450 10.3900 0.7450 10.3900 1.4600 10.4800 1.4600 10.4800 1.7000
                 10.3600 1.7000 10.3600 1.5800 10.2700 1.5800 10.2700 0.6000 9.7900 0.6000
                 9.7900 0.6200 9.1400 0.6200 9.1400 0.6000 7.6350 0.6000 7.6350 0.4800 7.5150 0.4800
                 7.5150 0.3600 7.7550 0.3600 7.7550 0.4800 8.6150 0.4800 8.6150 0.3800 8.8550 0.3800
                 8.8550 0.4800 9.2600 0.4800 9.2600 0.5000 9.6700 0.5000 9.6700 0.3800 9.9900 0.3800
                 9.9900 0.4800 10.4800 0.4800 ;
        POLYGON  10.1500 0.8400 10.0300 0.8400 10.0300 1.4600 9.9150 1.4600 9.9150 2.0200 9.7950 2.0200
                 9.7950 1.4600 9.1350 1.4600 9.1350 2.2000 8.4150 2.2000 8.4150 2.0100 7.0350 2.0100
                 7.0350 1.6600 6.7150 1.6600 6.7150 1.4400 6.3050 1.4400 6.3050 1.3200 6.8350 1.3200
                 6.8350 1.5400 7.1550 1.5400 7.1550 1.8900 8.5350 1.8900 8.5350 2.0800 9.0150 2.0800
                 9.0150 1.4600 8.6750 1.4600 8.6750 1.5300 8.5550 1.5300 8.5550 1.2900 8.6750 1.2900
                 8.6750 1.3400 9.0150 1.3400 9.0150 1.2800 9.2750 1.2800 9.2750 1.3400 9.9100 1.3400
                 9.9100 0.7200 10.1500 0.7200 ;
        POLYGON  9.0150 0.8400 8.8950 0.8400 8.8950 1.1700 8.4350 1.1700 8.4350 1.6500 8.7750 1.6500
                 8.7750 1.8400 8.8950 1.8400 8.8950 1.9600 8.6550 1.9600 8.6550 1.7700 8.3150 1.7700
                 8.3150 1.1700 7.1950 1.1700 7.1950 1.0500 8.7750 1.0500 8.7750 0.7200 9.0150 0.7200 ;
        POLYGON  8.1950 1.5600 7.9550 1.5600 7.9550 1.4200 7.3950 1.4200 7.3950 1.6500 7.5150 1.6500
                 7.5150 1.7700 7.2750 1.7700 7.2750 1.4200 6.9550 1.4200 6.9550 1.1400 6.1850 1.1400
                 6.1850 1.6600 5.8450 1.6600 5.8450 1.5400 6.0650 1.5400 6.0650 0.8600 5.9450 0.8600
                 5.9450 0.6200 6.0650 0.6200 6.0650 0.7400 6.1850 0.7400 6.1850 1.0200 6.9550 1.0200
                 6.9550 0.7800 7.0350 0.7800 7.0350 0.6600 7.1550 0.6600 7.1550 0.9000 7.0750 0.9000
                 7.0750 1.3000 8.0750 1.3000 8.0750 1.4400 8.1950 1.4400 ;
        POLYGON  7.6350 0.8400 7.3950 0.8400 7.3950 0.7200 7.2750 0.7200 7.2750 0.5400 6.8650 0.5400
                 6.8650 0.6600 6.7350 0.6600 6.7350 0.9000 6.6150 0.9000 6.6150 0.5400 6.7450 0.5400
                 6.7450 0.4200 7.3950 0.4200 7.3950 0.6000 7.5150 0.6000 7.5150 0.7200 7.6350 0.7200 ;
        POLYGON  6.6750 2.2300 6.4350 2.2300 6.4350 2.1400 5.9550 2.1400 5.9550 2.2000 4.8750 2.2000
                 4.8750 2.0600 4.3650 2.0600 4.3650 2.1300 4.3450 2.1300 4.3450 2.2500 4.2250 2.2500
                 4.2250 2.1300 2.6550 2.1300 2.6550 2.0850 2.2250 2.0850 2.2250 1.7250 2.2650 1.7250
                 2.2650 0.6100 2.3850 0.6100 2.3850 1.8450 2.3450 1.8450 2.3450 1.9650 2.7750 1.9650
                 2.7750 2.0100 4.2450 2.0100 4.2450 1.9400 4.9950 1.9400 4.9950 2.0800 5.8350 2.0800
                 5.8350 2.0200 6.5550 2.0200 6.5550 2.1100 6.6750 2.1100 ;
        POLYGON  5.9450 1.3400 5.7050 1.3400 5.7050 0.4800 5.2650 0.4800 5.2650 0.3600 5.8250 0.3600
                 5.8250 1.2200 5.9450 1.2200 ;
        POLYGON  5.5850 0.8600 5.4750 0.8600 5.4750 1.7200 5.3550 1.7200 5.3550 1.3400 3.4950 1.3400
                 3.4950 0.8800 3.0150 0.8800 3.0150 1.2400 3.0350 1.2400 3.0350 1.3600 2.7950 1.3600
                 2.7950 1.2400 2.8950 1.2400 2.8950 0.7600 3.6150 0.7600 3.6150 1.2200 5.3550 1.2200
                 5.3550 0.7400 5.4650 0.7400 5.4650 0.6200 5.5850 0.6200 ;
        POLYGON  5.1650 1.1000 4.2350 1.1000 4.2350 0.6200 4.3550 0.6200 4.3550 0.9800 5.0450 0.9800
                 5.0450 0.6200 5.1650 0.6200 ;
        POLYGON  5.1150 1.5800 3.8850 1.5800 3.8850 1.6500 3.6450 1.6500 3.6450 1.5300 3.7650 1.5300
                 3.7650 1.4600 5.1150 1.4600 ;
        POLYGON  4.7750 0.8600 4.6550 0.8600 4.6550 0.5000 4.1150 0.5000 4.1150 0.7200 3.9750 0.7200
                 3.9750 0.8000 3.7350 0.8000 3.7350 0.6800 3.8550 0.6800 3.8550 0.6000 3.9950 0.6000
                 3.9950 0.3800 4.7750 0.3800 ;
        POLYGON  3.8750 0.4800 3.7350 0.4800 3.7350 0.5600 2.7750 0.5600 2.7750 0.8600 2.6750 0.8600
                 2.6750 1.5200 2.8650 1.5200 2.8650 1.7600 2.7450 1.7600 2.7450 1.6400 2.5550 1.6400
                 2.5550 0.7400 2.6550 0.7400 2.6550 0.5600 2.5550 0.5600 2.5550 0.4900 2.1450 0.4900
                 2.1450 1.0900 1.7850 1.0900 1.7850 1.1100 1.5450 1.1100 1.5450 0.9700 2.0250 0.9700
                 2.0250 0.3700 2.6750 0.3700 2.6750 0.4400 3.6150 0.4400 3.6150 0.3600 3.8750 0.3600 ;
        POLYGON  1.0950 1.5800 0.9750 1.5800 0.9750 1.2000 0.3750 1.2000 0.3750 1.0800 0.9750 1.0800
                 0.9750 0.6800 1.0950 0.6800 ;
    END
END DFFNSRX1

MACRO DFFHQX8
    CLASS CORE ;
    FOREIGN DFFHQX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.5700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6550 0.6800 2.7750 2.1300 ;
        RECT  0.0700 1.0250 2.7750 1.1450 ;
        RECT  1.8150 0.6800 1.9350 2.1300 ;
        RECT  0.9750 0.6800 1.0950 2.1250 ;
        RECT  0.1350 0.6800 0.2550 2.1250 ;
        RECT  0.0700 0.8850 0.2550 1.1450 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.7700 1.0600 8.9200 1.4350 ;
        RECT  8.7250 1.0400 8.8450 1.4250 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.0400 1.0400 9.2150 1.4500 ;
        END
    END CK
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.5700 0.1800 ;
        RECT  8.8850 -0.1800 9.0050 0.6800 ;
        RECT  7.3250 0.4000 7.5650 0.5200 ;
        RECT  7.3250 -0.1800 7.4450 0.5200 ;
        RECT  5.4850 0.5000 5.7250 0.6200 ;
        RECT  5.4850 -0.1800 5.6050 0.6200 ;
        RECT  3.9150 -0.1800 4.0350 0.7300 ;
        RECT  3.0750 -0.1800 3.1950 0.7300 ;
        RECT  2.2350 -0.1800 2.3550 0.6700 ;
        RECT  1.3950 -0.1800 1.5150 0.6700 ;
        RECT  0.5550 -0.1800 0.6750 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.5700 2.7900 ;
        RECT  8.5850 1.8100 8.8250 1.9300 ;
        RECT  8.5850 1.8100 8.7050 2.7900 ;
        RECT  7.2450 2.0800 7.4850 2.2000 ;
        RECT  7.2450 2.0800 7.3650 2.7900 ;
        RECT  5.2650 2.2600 5.5050 2.7900 ;
        RECT  3.9150 2.0200 4.1550 2.1400 ;
        RECT  3.9150 2.0200 4.0350 2.7900 ;
        RECT  3.0750 1.4800 3.1950 2.7900 ;
        RECT  2.2350 1.3850 2.3550 2.7900 ;
        RECT  1.3950 1.3850 1.5150 2.7900 ;
        RECT  0.5550 1.3850 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.4250 0.8000 9.2450 0.8000 9.2450 0.9200 8.5250 0.9200 8.5250 1.5700 9.3250 1.5700
                 9.3250 1.8100 9.2050 1.8100 9.2050 1.6900 8.4650 1.6900 8.4650 2.2300 8.0450 2.2300
                 8.0450 2.2500 7.8050 2.2500 7.8050 2.2300 7.6450 2.2300 7.6450 1.9600 6.7050 1.9600
                 6.7050 2.2300 5.6250 2.2300 5.6250 2.1400 4.9450 2.1400 4.9450 2.0200 5.7450 2.0200
                 5.7450 2.1100 6.5850 2.1100 6.5850 1.2400 6.7450 1.2400 6.7450 1.1200 6.8650 1.1200
                 6.8650 1.3600 6.7050 1.3600 6.7050 1.8400 7.7650 1.8400 7.7650 2.1100 8.3450 2.1100
                 8.3450 1.5700 8.4050 1.5700 8.4050 0.8000 9.1250 0.8000 9.1250 0.6800 9.3050 0.6800
                 9.3050 0.4400 9.4250 0.4400 ;
        POLYGON  8.3050 0.6800 8.2850 0.6800 8.2850 1.3600 8.1250 1.3600 8.1250 1.9900 8.0050 1.9900
                 8.0050 1.3600 7.3450 1.3600 7.3450 1.3100 7.2250 1.3100 7.2250 1.1900 7.4650 1.1900
                 7.4650 1.2400 8.1650 1.2400 8.1650 0.5600 8.1850 0.5600 8.1850 0.4400 8.3050 0.4400 ;
        POLYGON  8.0450 1.1200 7.9250 1.1200 7.9250 0.7600 7.0850 0.7600 7.0850 0.4800 6.6050 0.4800
                 6.6050 1.1200 6.4050 1.1200 6.4050 0.8800 6.4850 0.8800 6.4850 0.4800 6.0050 0.4800
                 6.0050 0.8600 5.9850 0.8600 5.9850 1.5300 5.0250 1.5300 5.0250 1.6500 4.7850 1.6500
                 4.7850 1.5300 4.9050 1.5300 4.9050 1.4100 5.8650 1.4100 5.8650 0.8600 5.0650 0.8600
                 5.0650 0.5400 5.1850 0.5400 5.1850 0.7400 5.8850 0.7400 5.8850 0.3600 7.2050 0.3600
                 7.2050 0.6400 8.0450 0.6400 ;
        POLYGON  7.7850 1.0700 7.1050 1.0700 7.1050 1.6000 6.9450 1.6000 6.9450 1.7200 6.8250 1.7200
                 6.8250 1.4800 6.9850 1.4800 6.9850 1.0000 6.7250 1.0000 6.7250 0.6000 6.9650 0.6000
                 6.9650 0.8800 7.1050 0.8800 7.1050 0.9500 7.7850 0.9500 ;
        POLYGON  6.3650 0.7200 6.2450 0.7200 6.2450 1.9900 6.1250 1.9900 6.1250 1.9000 4.1550 1.9000
                 4.1550 1.3400 4.0350 1.3400 4.0350 1.2200 4.2750 1.2200 4.2750 1.7800 6.1250 1.7800
                 6.1250 0.6000 6.3650 0.6000 ;
        POLYGON  5.7250 1.1000 4.5150 1.1000 4.5150 1.5400 4.6350 1.5400 4.6350 1.6600 4.3950 1.6600
                 4.3950 1.1000 3.6150 1.1000 3.6150 2.1300 3.4950 2.1300 3.4950 1.1000 3.0550 1.1000
                 3.0550 1.2400 2.9350 1.2400 2.9350 0.9800 3.4950 0.9800 3.4950 0.6800 3.6150 0.6800
                 3.6150 0.9800 4.3350 0.9800 4.3350 0.6800 4.4550 0.6800 4.4550 0.8000 4.5150 0.8000
                 4.5150 0.9800 5.7250 0.9800 ;
    END
END DFFHQX8

MACRO DFFHQX4
    CLASS CORE ;
    FOREIGN DFFHQX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2100 1.3800 2.3300 2.0300 ;
        RECT  2.0300 1.3800 2.3300 1.5000 ;
        RECT  2.0300 0.6800 2.1500 1.5000 ;
        RECT  1.2300 1.0250 2.1500 1.1450 ;
        RECT  1.3700 1.0250 1.4900 2.0300 ;
        RECT  1.2300 0.7400 1.3800 1.1450 ;
        RECT  1.2600 1.0250 1.4900 1.2650 ;
        RECT  1.0100 0.7400 1.3800 0.8600 ;
        END
    END Q
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0400 0.5100 1.4450 ;
        RECT  0.3750 0.8450 0.4950 1.4450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.4050 1.2100 7.7500 1.3350 ;
        RECT  7.2650 1.2200 7.5250 1.3800 ;
        END
    END D
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.7100 -0.1800 7.8300 0.8300 ;
        RECT  5.7100 0.4900 5.9500 0.6100 ;
        RECT  5.8300 -0.1800 5.9500 0.6100 ;
        RECT  3.7100 0.4700 3.9500 0.5900 ;
        RECT  3.8300 -0.1800 3.9500 0.5900 ;
        RECT  2.5100 0.4700 2.7500 0.5900 ;
        RECT  2.5100 -0.1800 2.6300 0.5900 ;
        RECT  1.4900 -0.1800 1.7300 0.3200 ;
        RECT  0.5300 -0.1800 0.7700 0.3400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  7.3500 1.7400 7.4700 2.7900 ;
        RECT  5.6900 2.0100 5.8100 2.7900 ;
        RECT  3.6500 1.4700 3.7700 2.7900 ;
        RECT  2.6300 1.3800 2.7500 2.7900 ;
        RECT  1.7900 1.3800 1.9100 2.7900 ;
        RECT  0.9500 1.3800 1.0700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.3500 1.6200 8.2500 1.6200 8.2500 1.6500 8.0100 1.6500 8.0100 1.6200 7.0300 1.6200
                 7.0300 2.2300 6.1150 2.2300 6.1150 1.8900 4.9900 1.8900 4.9900 2.2500 4.0900 2.2500
                 4.0900 2.1300 4.8700 2.1300 4.8700 0.9700 5.1100 0.9700 5.1100 1.0900 4.9900 1.0900
                 4.9900 1.7700 6.2350 1.7700 6.2350 2.1100 6.9100 2.1100 6.9100 1.3300 6.7900 1.3300
                 6.7900 1.2100 7.0300 1.2100 7.0300 1.5000 8.2300 1.5000 8.2300 0.8500 8.1300 0.8500
                 8.1300 0.5900 8.2500 0.5900 8.2500 0.7300 8.3500 0.7300 ;
        POLYGON  8.1100 1.0900 7.1500 1.0900 7.1500 0.9700 7.2900 0.9700 7.2900 0.5300 6.4300 0.5300
                 6.4300 0.8500 6.3850 0.8500 6.3850 1.2100 6.4300 1.2100 6.4300 1.3300 6.1900 1.3300
                 6.1900 1.2100 6.2650 1.2100 6.2650 0.8500 5.4700 0.8500 5.4700 0.5300 4.3900 0.5300
                 4.3900 0.9700 4.5100 0.9700 4.5100 1.0900 4.2700 1.0900 4.2700 0.8300 3.4700 0.8300
                 3.4700 0.5300 2.9900 0.5300 2.9900 0.8300 2.2700 0.8300 2.2700 0.5600 1.8450 0.5600
                 1.8450 0.6200 0.7850 0.6200 0.7850 0.6800 0.2550 0.6800 0.2550 0.9200 0.2400 0.9200
                 0.2400 1.5650 0.5500 1.5650 0.5500 1.8050 0.4300 1.8050 0.4300 1.6850 0.1200 1.6850
                 0.1200 0.8000 0.1350 0.8000 0.1350 0.5600 0.6650 0.5600 0.6650 0.5000 1.7250 0.5000
                 1.7250 0.4400 2.3900 0.4400 2.3900 0.7100 2.8700 0.7100 2.8700 0.4100 3.5900 0.4100
                 3.5900 0.7100 4.2700 0.7100 4.2700 0.4100 5.5900 0.4100 5.5900 0.7300 6.3100 0.7300
                 6.3100 0.4100 7.4100 0.4100 7.4100 0.9700 8.1100 0.9700 ;
        POLYGON  7.1700 0.7700 6.6700 0.7700 6.6700 1.9900 6.5500 1.9900 6.5500 1.5700 5.9500 1.5700
                 5.9500 1.3500 5.5900 1.3500 5.5900 1.3300 5.4700 1.3300 5.4700 1.2100 5.7100 1.2100
                 5.7100 1.2300 6.0700 1.2300 6.0700 1.4500 6.5500 1.4500 6.5500 0.6500 7.1700 0.6500 ;
        POLYGON  6.0700 1.1100 5.8300 1.1100 5.8300 1.0900 5.3500 1.0900 5.3500 1.6500 5.1100 1.6500
                 5.1100 1.5300 5.2300 1.5300 5.2300 0.7700 5.1100 0.7700 5.1100 0.6500 5.3500 0.6500
                 5.3500 0.9700 5.9500 0.9700 5.9500 0.9900 6.0700 0.9900 ;
        POLYGON  4.7900 0.7700 4.7500 0.7700 4.7500 1.3300 4.4100 1.3300 4.4100 1.9900 4.2900 1.9900
                 4.2900 1.3300 3.3700 1.3300 3.3700 1.1900 3.6100 1.1900 3.6100 1.2100 4.6300 1.2100
                 4.6300 0.7700 4.5500 0.7700 4.5500 0.6500 4.7900 0.6500 ;
        POLYGON  3.9700 1.0900 3.7300 1.0900 3.7300 1.0700 3.2500 1.0700 3.2500 1.4500 3.2900 1.4500
                 3.2900 1.9900 3.1700 1.9900 3.1700 1.5700 3.1300 1.5700 3.1300 1.0700 2.4100 1.0700
                 2.4100 1.2600 2.2900 1.2600 2.2900 0.9500 3.1100 0.9500 3.1100 0.6500 3.3500 0.6500
                 3.3500 0.7700 3.2300 0.7700 3.2300 0.9500 3.8500 0.9500 3.8500 0.9700 3.9700 0.9700 ;
    END
END DFFHQX4

MACRO DFFHQX2
    CLASS CORE ;
    FOREIGN DFFHQX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2850 1.0000 0.4050 1.2400 ;
        RECT  0.0700 1.0000 0.4050 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.1200 1.7550 1.3550 ;
        RECT  1.1750 1.1200 1.4350 1.3800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5150 0.6400 5.6350 1.1800 ;
        RECT  5.4550 1.0600 5.5750 2.2100 ;
        RECT  5.2900 1.1750 5.5750 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  5.9950 -0.1800 6.1150 0.7800 ;
        RECT  4.9150 0.5800 5.1550 0.7000 ;
        RECT  4.9150 -0.1800 5.0350 0.7000 ;
        RECT  3.0150 0.5800 3.2550 0.7000 ;
        RECT  3.0150 -0.1800 3.1350 0.7000 ;
        RECT  1.4950 0.6000 1.7350 0.7200 ;
        RECT  1.6150 -0.1800 1.7350 0.7200 ;
        RECT  0.1350 -0.1800 0.2550 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  5.8750 1.5600 5.9950 2.7900 ;
        RECT  5.0350 1.5600 5.1550 2.7900 ;
        RECT  3.2150 2.2300 3.4550 2.7900 ;
        RECT  1.4150 1.7600 1.5350 2.7900 ;
        RECT  0.1450 1.4600 0.2650 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.5350 1.4400 6.4750 1.4400 6.4750 2.0800 6.3550 2.0800 6.3550 1.4400 5.7550 1.4400
                 5.7550 1.2000 5.8750 1.2000 5.8750 1.3200 6.4150 1.3200 6.4150 0.6400 6.5350 0.6400 ;
        POLYGON  6.2350 1.2000 6.1150 1.2000 6.1150 1.0200 5.7550 1.0200 5.7550 0.5200 5.3950 0.5200
                 5.3950 0.9400 4.8950 0.9400 4.8950 1.4200 4.6150 1.4200 4.6150 1.8100 4.4550 1.8100
                 4.4550 2.2100 4.3350 2.2100 4.3350 1.6900 4.4950 1.6900 4.4950 1.3000 4.7750 1.3000
                 4.7750 0.9400 4.6600 0.9400 4.6600 0.8000 4.2750 0.8000 4.2750 0.6800 4.7800 0.6800
                 4.7800 0.8200 5.2750 0.8200 5.2750 0.4000 5.8750 0.4000 5.8750 0.9000 6.2350 0.9000 ;
        POLYGON  4.6550 1.1800 3.9750 1.1800 3.9750 1.6100 3.8550 1.6100 3.8550 1.0600 3.8750 1.0600
                 3.8750 0.5000 3.4950 0.5000 3.4950 0.9400 2.8550 0.9400 2.8550 1.5900 2.7350 1.5900
                 2.7350 0.5600 2.0150 0.5600 2.0150 0.9600 2.0350 0.9600 2.0350 1.4000 1.9150 1.4000
                 1.9150 1.0800 1.8950 1.0800 1.8950 0.9600 1.2550 0.9600 1.2550 0.5600 0.6850 0.5600
                 0.6850 1.5800 0.5650 1.5800 0.5650 0.4400 1.1550 0.4400 1.1550 0.3600 1.3950 0.3600
                 1.3950 0.4800 1.3750 0.4800 1.3750 0.8400 1.8950 0.8400 1.8950 0.4400 2.8550 0.4400
                 2.8550 0.8200 3.3750 0.8200 3.3750 0.3800 3.9950 0.3800 3.9950 1.0600 4.6550 1.0600 ;
        POLYGON  4.3750 1.5700 4.2150 1.5700 4.2150 2.1100 2.9050 2.1100 2.9050 2.2500 2.2550 2.2500
                 2.2550 1.6400 1.0550 1.6400 1.0550 2.0900 0.9350 2.0900 0.9350 0.8000 0.8950 0.8000
                 0.8950 0.6800 1.1350 0.6800 1.1350 0.8000 1.0550 0.8000 1.0550 1.5200 2.2550 1.5200
                 2.2550 1.3500 2.3750 1.3500 2.3750 2.1300 2.7850 2.1300 2.7850 1.9900 4.0950 1.9900
                 4.0950 1.4500 4.2550 1.4500 4.2550 1.3300 4.3750 1.3300 ;
        POLYGON  3.9350 1.8700 3.6150 1.8700 3.6150 1.1900 3.0150 1.1900 3.0150 1.0700 3.6150 1.0700
                 3.6150 0.7400 3.6350 0.7400 3.6350 0.6200 3.7550 0.6200 3.7550 0.8600 3.7350 0.8600
                 3.7350 1.7500 3.9350 1.7500 ;
        POLYGON  3.4950 1.8300 2.6150 1.8300 2.6150 2.0100 2.4950 2.0100 2.4950 0.8000 2.1350 0.8000
                 2.1350 0.6800 2.6150 0.6800 2.6150 1.7100 3.3750 1.7100 3.3750 1.3500 3.4950 1.3500 ;
    END
END DFFHQX2

MACRO DFFHQX1
    CLASS CORE ;
    FOREIGN DFFHQX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CK
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7500 1.0900 0.8700 1.4550 ;
        RECT  0.6500 1.0900 0.8700 1.4500 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.1950 1.2050 5.4950 1.4200 ;
        RECT  5.2350 1.1800 5.4950 1.4200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1450 1.2950 0.2650 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4350 ;
        END
    END Q
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.3950 0.4500 5.6350 0.5700 ;
        RECT  5.3950 -0.1800 5.5150 0.5700 ;
        RECT  3.7950 0.4100 4.0350 0.5300 ;
        RECT  3.9150 -0.1800 4.0350 0.5300 ;
        RECT  2.0150 -0.1800 2.1350 0.6800 ;
        RECT  0.5550 -0.1800 0.6750 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.3950 1.5400 5.5150 2.7900 ;
        RECT  3.7950 2.0900 4.0350 2.2100 ;
        RECT  3.7950 2.0900 3.9150 2.7900 ;
        RECT  1.7150 2.0100 1.9550 2.1300 ;
        RECT  1.7150 2.0100 1.8350 2.7900 ;
        RECT  0.5650 1.8500 0.6850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.0550 0.7800 6.0350 0.7800 6.0350 1.3000 5.9950 1.3000 5.9950 1.7100 5.8750 1.7100
                 5.8750 1.1800 5.9150 1.1800 5.9150 0.8100 5.0150 0.8100 5.0150 0.4800 4.5350 0.4800
                 4.5350 1.1000 4.4150 1.1000 4.4150 0.7700 3.5550 0.7700 3.5550 0.4800 3.0750 0.4800
                 3.0750 0.9800 3.0350 0.9800 3.0350 1.1000 3.0150 1.1000 3.0150 1.1600 2.4550 1.1600
                 2.4550 1.3900 2.3350 1.3900 2.3350 1.0400 2.8950 1.0400 2.8950 0.8600 2.9550 0.8600
                 2.9550 0.3600 3.6750 0.3600 3.6750 0.6500 4.4150 0.6500 4.4150 0.3600 5.1350 0.3600
                 5.1350 0.6900 5.8100 0.6900 5.8100 0.6600 5.9350 0.6600 5.9350 0.5400 6.0550 0.5400 ;
        POLYGON  5.7950 1.0600 5.0150 1.0600 5.0150 1.9700 4.4750 1.9700 4.4750 2.1300 4.5950 2.1300
                 4.5950 2.2500 4.3550 2.2500 4.3550 1.9700 3.2550 1.9700 3.2550 2.2300 2.0750 2.2300
                 2.0750 1.8900 1.4000 1.8900 1.4000 1.9800 1.1050 1.9800 1.1050 2.1000 0.9850 2.1000
                 0.9850 1.8600 0.9950 1.8600 0.9950 1.2900 1.0350 1.2900 1.0350 0.6800 1.1550 0.6800
                 1.1550 1.4100 1.1150 1.4100 1.1150 1.8600 1.2800 1.8600 1.2800 1.7700 2.1950 1.7700
                 2.1950 2.1100 3.1350 2.1100 3.1350 1.2500 3.2750 1.2500 3.2750 1.1300 3.3950 1.1300
                 3.3950 1.3700 3.2550 1.3700 3.2550 1.8500 4.8950 1.8500 4.8950 0.9300 5.0150 0.9300
                 5.0150 0.9400 5.7950 0.9400 ;
        POLYGON  4.8950 0.7200 4.7750 0.7200 4.7750 1.3400 4.6750 1.3400 4.6750 1.7300 4.5550 1.7300
                 4.5550 1.3700 3.7550 1.3700 3.7550 1.1300 3.8750 1.1300 3.8750 1.2500 4.5550 1.2500
                 4.5550 1.2200 4.6550 1.2200 4.6550 0.6000 4.8950 0.6000 ;
        POLYGON  4.1950 1.1300 4.0750 1.1300 4.0750 1.0100 3.6350 1.0100 3.6350 1.6100 3.4950 1.6100
                 3.4950 1.7300 3.3750 1.7300 3.3750 1.4900 3.5150 1.4900 3.5150 1.0100 3.1950 1.0100
                 3.1950 0.6000 3.4350 0.6000 3.4350 0.8900 4.1950 0.8900 ;
        POLYGON  2.8350 0.7200 2.3750 0.7200 2.3750 0.9200 2.2150 0.9200 2.2150 1.5100 2.5750 1.5100
                 2.5750 1.4700 2.6950 1.4700 2.6950 1.9900 2.5750 1.9900 2.5750 1.6300 1.5950 1.6300
                 1.5950 1.3700 1.5150 1.3700 1.5150 1.1300 1.7150 1.1300 1.7150 1.5100 2.0950 1.5100
                 2.0950 0.8000 2.2550 0.8000 2.2550 0.6000 2.8350 0.6000 ;
        POLYGON  1.9750 1.3900 1.8550 1.3900 1.8550 1.0100 1.3950 1.0100 1.3950 1.5300 1.4750 1.5300
                 1.4750 1.6500 1.2350 1.6500 1.2350 1.5300 1.2750 1.5300 1.2750 0.5600 0.9150 0.5600
                 0.9150 0.9700 0.5300 0.9700 0.5300 1.2400 0.4100 1.2400 0.4100 0.8500 0.7950 0.8500
                 0.7950 0.4400 1.7150 0.4400 1.7150 0.8900 1.9750 0.8900 ;
    END
END DFFHQX1

MACRO CLKXOR2X8
    CLASS CORE ;
    FOREIGN CLKXOR2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3650 0.9600 3.4850 1.3600 ;
        RECT  3.2050 0.9400 3.4650 1.1650 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2550 1.1100 5.4950 1.2300 ;
        RECT  5.2900 1.1100 5.4400 1.4350 ;
        RECT  4.6750 1.0400 5.4100 1.1600 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7250 1.4100 2.8450 2.2100 ;
        RECT  2.5950 0.7150 2.8350 0.8350 ;
        RECT  2.5450 1.4100 2.8450 1.5300 ;
        RECT  0.1350 0.7600 2.7150 0.8800 ;
        RECT  0.3600 1.2900 2.6650 1.4100 ;
        RECT  1.8850 1.2900 2.0050 2.2100 ;
        RECT  1.7550 0.7100 1.9950 0.8800 ;
        RECT  1.0450 1.2900 1.1650 2.2100 ;
        RECT  0.9150 0.7100 1.1550 0.8800 ;
        RECT  0.3600 0.7600 0.5100 1.1450 ;
        RECT  0.2050 1.4100 0.4800 1.5300 ;
        RECT  0.3600 0.7600 0.4800 1.5300 ;
        RECT  0.2050 1.4100 0.3250 2.2100 ;
        RECT  0.1350 0.6400 0.2550 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.2350 -0.1800 5.3550 0.6800 ;
        RECT  3.0150 0.4600 3.2550 0.5800 ;
        RECT  3.0150 -0.1800 3.1350 0.5800 ;
        RECT  2.2350 -0.1800 2.3550 0.6400 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  4.9750 1.7600 5.0950 2.7900 ;
        RECT  3.0850 2.0000 3.3250 2.1500 ;
        RECT  3.0850 2.0000 3.2050 2.7900 ;
        RECT  2.3050 1.5300 2.4250 2.7900 ;
        RECT  1.4650 1.5300 1.5850 2.7900 ;
        RECT  0.6250 1.5300 0.7450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7750 0.9200 5.7350 0.9200 5.7350 1.6750 5.5750 1.6750 5.5750 1.9300 5.4550 1.9300
                 5.4550 1.5550 5.6150 1.5550 5.6150 0.9200 4.4550 0.9200 4.4550 1.2800 4.5750 1.2800
                 4.5750 1.4000 4.3350 1.4000 4.3350 1.0400 3.9750 1.0400 3.9750 1.1200 3.8550 1.1200
                 3.8550 0.8800 3.9750 0.8800 3.9750 0.9200 4.3350 0.9200 4.3350 0.8000 5.6150 0.8000
                 5.6150 0.5600 5.6550 0.5600 5.6550 0.4400 5.7750 0.4400 ;
        POLYGON  5.0750 1.6400 4.0350 1.6400 4.0350 2.0100 3.9150 2.0100 3.9150 1.6400 3.6150 1.6400
                 3.6150 0.6000 3.8750 0.6000 3.8750 0.7200 3.7350 0.7200 3.7350 1.5200 4.9550 1.5200
                 4.9550 1.3700 5.0750 1.3700 ;
        POLYGON  4.4550 2.2100 4.3600 2.2100 4.3600 2.2500 3.4450 2.2500 3.4450 1.8800 3.1800 1.8800
                 3.1800 1.7600 2.9650 1.7600 2.9650 1.1700 1.9350 1.1700 1.9350 1.0500 2.9650 1.0500
                 2.9650 0.7000 3.3750 0.7000 3.3750 0.3600 4.2350 0.3600 4.2350 0.6800 4.1150 0.6800
                 4.1150 0.4800 3.4950 0.4800 3.4950 0.8200 3.0850 0.8200 3.0850 1.6400 3.3000 1.6400
                 3.3000 1.7600 3.5650 1.7600 3.5650 2.1300 4.2400 2.1300 4.2400 2.0900 4.3350 2.0900
                 4.3350 1.7600 4.4550 1.7600 ;
    END
END CLKXOR2X8

MACRO CLKXOR2X4
    CLASS CORE ;
    FOREIGN CLKXOR2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.1800 2.1750 1.3450 ;
        RECT  1.7550 1.1800 2.0150 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8400 1.1750 3.9900 1.4350 ;
        RECT  3.8400 1.0400 3.9600 1.4350 ;
        RECT  3.1150 1.0400 3.9600 1.1600 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 1.7400 1.5750 2.2100 ;
        RECT  1.2150 0.7000 1.5150 0.8200 ;
        RECT  1.3950 0.5800 1.5150 0.8200 ;
        RECT  1.2750 1.7400 1.5750 1.8600 ;
        RECT  1.2750 1.3200 1.3950 1.8600 ;
        RECT  0.6500 0.8400 1.3350 0.9600 ;
        RECT  1.2150 0.7000 1.3350 0.9600 ;
        RECT  0.6500 1.3200 1.3950 1.4400 ;
        RECT  0.6500 1.1750 0.8000 1.4400 ;
        RECT  0.6500 0.7900 0.7700 1.5600 ;
        RECT  0.6150 1.4400 0.7350 2.2100 ;
        RECT  0.5550 0.6700 0.6750 0.9100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.6750 -0.1800 3.7950 0.6800 ;
        RECT  1.8150 -0.1800 1.9350 0.7200 ;
        RECT  0.9750 -0.1800 1.0950 0.7200 ;
        RECT  0.1350 -0.1800 0.2550 0.7200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.6750 1.8400 3.7950 2.7900 ;
        RECT  1.8750 2.0800 2.1150 2.2000 ;
        RECT  1.8750 2.0800 1.9950 2.7900 ;
        RECT  1.0350 1.5600 1.1550 2.7900 ;
        RECT  0.1950 1.5600 0.3150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.2300 1.9600 4.2150 1.9600 4.2150 2.0800 4.0950 2.0800 4.0950 1.8400 4.1100 1.8400
                 4.1100 0.9200 2.9950 0.9200 2.9950 1.3600 3.3550 1.3600 3.3550 1.4800 2.8750 1.4800
                 2.8750 1.1000 2.5350 1.1000 2.5350 0.8600 2.6550 0.8600 2.6550 0.9800 2.8750 0.9800
                 2.8750 0.8000 4.0950 0.8000 4.0950 0.4400 4.2150 0.4400 4.2150 0.5600 4.2300 0.5600 ;
        POLYGON  3.6350 1.7200 2.7350 1.7200 2.7350 2.0100 2.6150 2.0100 2.6150 1.7200 2.2950 1.7200
                 2.2950 0.6000 2.7550 0.6000 2.7550 0.7200 2.4150 0.7200 2.4150 1.6000 3.5150 1.6000
                 3.5150 1.3400 3.6350 1.3400 ;
        POLYGON  3.1550 2.2500 2.2350 2.2500 2.2350 1.9600 1.9700 1.9600 1.9700 1.6200 1.5150 1.6200
                 1.5150 1.2000 1.2550 1.2000 1.2550 1.0800 1.5150 1.0800 1.5150 0.9400 2.0550 0.9400
                 2.0550 0.3600 3.1150 0.3600 3.1150 0.6800 2.9950 0.6800 2.9950 0.4800 2.1750 0.4800
                 2.1750 1.0600 1.6350 1.0600 1.6350 1.5000 2.0900 1.5000 2.0900 1.8400 2.3550 1.8400
                 2.3550 2.1300 3.0350 2.1300 3.0350 1.8400 3.1550 1.8400 ;
    END
END CLKXOR2X4

MACRO CLKXOR2X2
    CLASS CORE ;
    FOREIGN CLKXOR2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 1.2200 1.3350 1.4600 ;
        RECT  0.8850 1.2300 1.3350 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8150 1.1800 3.1750 1.3000 ;
        RECT  2.3350 1.1800 2.5950 1.3800 ;
        RECT  2.2550 1.1400 2.4950 1.3000 ;
        RECT  1.6950 1.3400 1.9350 1.4600 ;
        RECT  1.8150 1.1800 1.9350 1.4600 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5950 1.7400 0.7150 2.2100 ;
        RECT  0.4050 0.7400 0.6750 0.8600 ;
        RECT  0.5550 0.6200 0.6750 0.8600 ;
        RECT  0.4050 1.7400 0.7150 1.8600 ;
        RECT  0.4050 0.7400 0.5250 1.8600 ;
        RECT  0.3600 0.8850 0.5250 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.7350 -0.1800 2.8550 0.7800 ;
        RECT  0.9750 -0.1800 1.0950 0.7300 ;
        RECT  0.1350 -0.1800 0.2550 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.6150 1.7400 2.7350 2.7900 ;
        RECT  1.0150 2.2200 1.2550 2.7900 ;
        RECT  0.1650 1.5600 0.2850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.4150 1.7400 3.1550 1.7400 3.1550 1.8600 3.0350 1.8600 3.0350 1.6200 2.3350 1.6200
                 2.3350 2.2400 2.0550 2.2400 2.0550 2.1200 2.2150 2.1200 2.2150 1.5000 3.1550 1.5000
                 3.1550 1.6200 3.2950 1.6200 3.2950 0.7800 3.1550 0.7800 3.1550 0.5400 3.2750 0.5400
                 3.2750 0.6600 3.4150 0.6600 ;
        POLYGON  2.8550 1.0600 2.6150 1.0600 2.6150 1.0200 1.5750 1.0200 1.5750 1.5800 1.6750 1.5800
                 1.6750 1.8600 1.5550 1.8600 1.5550 1.7000 1.4550 1.7000 1.4550 0.6000 1.6950 0.6000
                 1.6950 0.7200 1.5750 0.7200 1.5750 0.9000 2.7350 0.9000 2.7350 0.9400 2.8550 0.9400 ;
        POLYGON  2.2150 0.7800 2.0950 0.7800 2.0950 0.4800 1.3350 0.4800 1.3350 1.1000 0.7650 1.1000
                 0.7650 1.5000 0.9550 1.5000 0.9550 1.5800 1.1400 1.5800 1.1400 1.9800 1.8150 1.9800
                 1.8150 1.8600 1.9750 1.8600 1.9750 1.7400 2.0950 1.7400 2.0950 1.9800 1.9350 1.9800
                 1.9350 2.1000 1.0200 2.1000 1.0200 1.7000 0.8350 1.7000 0.8350 1.6200 0.6450 1.6200
                 0.6450 0.9800 1.2150 0.9800 1.2150 0.3600 2.2150 0.3600 ;
    END
END CLKXOR2X2

MACRO CLKXOR2X1
    CLASS CORE ;
    FOREIGN CLKXOR2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8550 1.2800 0.9750 1.5600 ;
        RECT  0.6800 1.4400 0.9750 1.5600 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4550 1.1800 2.8350 1.3000 ;
        RECT  2.0450 1.1800 2.3050 1.3800 ;
        RECT  1.9150 1.1400 2.1550 1.3000 ;
        RECT  1.3350 1.3600 1.5750 1.4800 ;
        RECT  1.4550 1.1800 1.5750 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 1.2950 0.2900 2.2100 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        RECT  0.1350 0.6800 0.2550 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.3950 -0.1800 2.5150 0.7800 ;
        RECT  0.4950 0.5500 0.7350 0.6700 ;
        RECT  0.6150 -0.1800 0.7350 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.2750 1.7400 2.3950 2.7900 ;
        RECT  0.5900 2.1600 0.8300 2.2800 ;
        RECT  0.5900 2.1600 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0750 1.7400 2.8150 1.7400 2.8150 1.8600 2.6950 1.8600 2.6950 1.6200 1.9550 1.6200
                 1.9550 2.2400 1.7150 2.2400 1.7150 2.1200 1.8350 2.1200 1.8350 1.5000 2.8150 1.5000
                 2.8150 1.6200 2.9550 1.6200 2.9550 0.7800 2.8150 0.7800 2.8150 0.5400 2.9350 0.5400
                 2.9350 0.6600 3.0750 0.6600 ;
        POLYGON  2.5150 1.0600 2.2750 1.0600 2.2750 1.0200 1.2150 1.0200 1.2150 1.6800 1.3100 1.6800
                 1.3100 1.8000 1.0700 1.8000 1.0700 1.6800 1.0950 1.6800 1.0950 0.6000 1.3350 0.6000
                 1.3350 0.7200 1.2150 0.7200 1.2150 0.9000 2.3950 0.9000 2.3950 0.9400 2.5150 0.9400 ;
        POLYGON  1.8750 0.7800 1.7550 0.7800 1.7550 0.4800 0.9750 0.4800 0.9750 1.1600 0.5500 1.1600
                 0.5500 1.2800 0.5300 1.2800 0.5300 1.9200 1.4750 1.9200 1.4750 1.8600 1.5500 1.8600
                 1.5500 1.7400 1.6700 1.7400 1.6700 1.9800 1.5950 1.9800 1.5950 2.0400 0.4100 2.0400
                 0.4100 1.0400 0.8550 1.0400 0.8550 0.3600 1.8750 0.3600 ;
    END
END CLKXOR2X1

MACRO CLKMX2X8
    CLASS CORE ;
    FOREIGN CLKMX2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.8000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 1.1200 1.5050 1.2400 ;
        RECT  0.6450 1.5000 1.3850 1.6200 ;
        RECT  1.2650 1.1200 1.3850 1.6200 ;
        RECT  0.6450 1.1750 0.7650 1.6200 ;
        RECT  0.3600 1.1750 0.7650 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1100 1.1450 1.3800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0800 2.5400 1.4600 ;
        RECT  2.2800 1.0800 2.5400 1.2750 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7250 0.7650 5.4650 0.8850 ;
        RECT  5.3450 0.6450 5.4650 0.8850 ;
        RECT  5.3400 0.7650 5.4600 2.2050 ;
        RECT  2.9700 1.2250 5.4600 1.3450 ;
        RECT  4.4450 0.7150 4.6850 0.8850 ;
        RECT  4.5000 1.2250 4.6200 2.2050 ;
        RECT  3.6050 0.7150 3.8450 0.8350 ;
        RECT  3.6600 1.2250 3.7800 2.2100 ;
        RECT  2.9700 1.1750 3.1200 1.4350 ;
        RECT  2.8200 1.3450 3.0900 1.4650 ;
        RECT  2.9700 0.6000 3.0900 1.4650 ;
        RECT  2.7650 0.6000 3.0900 0.7200 ;
        RECT  2.8200 1.3450 2.9400 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.8000 0.1800 ;
        RECT  4.9250 -0.1800 5.0450 0.6450 ;
        RECT  4.0850 -0.1800 4.2050 0.6450 ;
        RECT  3.2450 -0.1800 3.3650 0.6450 ;
        RECT  2.3450 0.4600 2.5850 0.5800 ;
        RECT  2.3450 -0.1800 2.4650 0.5800 ;
        RECT  0.8250 -0.1800 0.9450 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.8000 2.7900 ;
        RECT  4.9200 1.4650 5.0400 2.7900 ;
        RECT  4.0800 1.4650 4.2000 2.7900 ;
        RECT  3.2400 1.4650 3.3600 2.7900 ;
        RECT  2.4000 1.5800 2.5200 2.7900 ;
        RECT  0.9600 1.7400 1.2000 2.1400 ;
        RECT  0.9600 1.7400 1.0800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.8000 1.2150 2.6800 1.2150 2.6800 0.9600 2.1600 0.9600 2.1600 1.7800 1.7800 1.7800
                 1.7800 2.2000 1.6600 2.2000 1.6600 1.6600 2.0400 1.6600 2.0400 0.9600 1.9850 0.9600
                 1.9850 0.7500 1.7650 0.7500 1.7650 0.5000 1.8850 0.5000 1.8850 0.6300 2.1050 0.6300
                 2.1050 0.8400 2.8000 0.8400 ;
        POLYGON  1.9200 1.5400 1.6250 1.5400 1.6250 0.9900 0.2400 0.9900 0.2400 1.5550 0.5250 1.5550
                 0.5250 1.9200 0.4050 1.9200 0.4050 1.6750 0.1200 1.6750 0.1200 0.7500 0.3450 0.7500
                 0.3450 0.5000 0.4650 0.5000 0.4650 0.8700 1.7450 0.8700 1.7450 0.8800 1.8650 0.8800
                 1.8650 1.0000 1.7450 1.0000 1.7450 1.4200 1.9200 1.4200 ;
    END
END CLKMX2X8

MACRO CLKMX2X6
    CLASS CORE ;
    FOREIGN CLKMX2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4100 1.5550 1.1700 1.6750 ;
        RECT  1.0500 1.3500 1.1700 1.6750 ;
        RECT  0.4100 1.1950 0.5300 1.6750 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0450 0.8500 1.4350 ;
        RECT  0.7300 1.0350 0.8500 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8700 1.2150 2.2500 1.4350 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.8700 1.2150 1.9900 1.4550 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2100 1.4300 4.3300 2.2100 ;
        RECT  3.9900 0.8000 4.2900 0.9200 ;
        RECT  4.1700 0.4050 4.2900 0.9200 ;
        RECT  4.0300 1.4300 4.3300 1.5500 ;
        RECT  4.0300 1.1900 4.1500 1.5500 ;
        RECT  3.3300 1.0400 4.1100 1.3100 ;
        RECT  3.9900 0.8000 4.1100 1.3100 ;
        RECT  3.3700 1.0400 3.4900 2.2100 ;
        RECT  3.3300 0.4050 3.4500 1.3100 ;
        RECT  2.6700 1.1900 4.1500 1.3100 ;
        RECT  2.6700 1.1750 2.8300 1.4350 ;
        RECT  2.5300 1.3600 2.7900 1.4800 ;
        RECT  2.6700 0.6300 2.7900 1.4800 ;
        RECT  2.4300 0.6300 2.7900 0.7500 ;
        RECT  2.5300 1.3600 2.6500 2.2100 ;
        RECT  2.4300 0.4000 2.5500 0.7500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  3.7500 -0.1800 3.8700 0.9200 ;
        RECT  2.9100 -0.1800 3.0300 0.9200 ;
        RECT  2.0100 -0.1800 2.1300 0.7400 ;
        RECT  0.7300 -0.1800 0.8500 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  3.7900 1.4300 3.9100 2.7900 ;
        RECT  2.9500 1.4300 3.0700 2.7900 ;
        RECT  2.1100 1.5550 2.2300 2.7900 ;
        RECT  0.5700 1.7950 0.6900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4900 1.2400 2.3700 1.2400 2.3700 0.9900 1.7500 0.9900 1.7500 1.8400 1.4300 1.8400
                 1.4300 2.2100 1.3100 2.2100 1.3100 1.7200 1.6300 1.7200 1.6300 0.9900 1.4700 0.9900
                 1.4700 0.6750 1.3700 0.6750 1.3700 0.4350 1.4900 0.4350 1.4900 0.5550 1.5900 0.5550
                 1.5900 0.8700 2.4900 0.8700 ;
        POLYGON  1.5100 1.6000 1.3900 1.6000 1.3900 1.2300 1.2300 1.2300 1.2300 0.9150 0.2400 0.9150
                 0.2400 1.5550 0.2700 1.5550 0.2700 2.0350 0.1500 2.0350 0.1500 1.6750 0.1200 1.6750
                 0.1200 0.6750 0.2500 0.6750 0.2500 0.5000 0.3700 0.5000 0.3700 0.7950 1.3500 0.7950
                 1.3500 1.1100 1.5100 1.1100 ;
    END
END CLKMX2X6

MACRO CLKMX2X4
    CLASS CORE ;
    FOREIGN CLKMX2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.0600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1460  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9200 1.2000 1.2000 1.3200 ;
        RECT  0.3600 1.6000 1.0400 1.7200 ;
        RECT  0.9200 1.2000 1.0400 1.7200 ;
        RECT  0.3600 1.1750 0.5100 1.7200 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0250 0.8000 1.4800 ;
        RECT  0.6800 1.0000 0.8000 1.4800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.2300 2.3300 1.3950 ;
        RECT  1.8600 1.2750 2.1900 1.4050 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2400 1.4400 3.3600 2.2100 ;
        RECT  3.2200 0.5900 3.3400 0.8300 ;
        RECT  3.0600 1.4400 3.3600 1.5600 ;
        RECT  3.0400 0.7100 3.3400 0.8300 ;
        RECT  2.5600 1.3200 3.1800 1.4400 ;
        RECT  2.5600 0.7600 3.1600 0.8800 ;
        RECT  2.5600 1.1750 2.8300 1.4400 ;
        RECT  2.4000 1.5150 2.6800 1.6350 ;
        RECT  2.5600 0.6500 2.6800 1.6350 ;
        RECT  2.3200 0.6500 2.6800 0.7700 ;
        RECT  2.4000 1.5150 2.5200 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.0600 0.1800 ;
        RECT  3.6400 -0.1800 3.7600 0.6400 ;
        RECT  2.8000 -0.1800 2.9200 0.6400 ;
        RECT  1.9000 0.4600 2.1400 0.5800 ;
        RECT  1.9000 -0.1800 2.0200 0.5800 ;
        RECT  0.6800 -0.1800 0.8000 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.0600 2.7900 ;
        RECT  3.6600 1.5600 3.7800 2.7900 ;
        RECT  2.8200 1.5600 2.9400 2.7900 ;
        RECT  1.9800 1.5600 2.1000 2.7900 ;
        RECT  0.6400 1.8400 0.7600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4400 1.1100 1.7400 1.1100 1.7400 1.8400 1.4000 1.8400 1.4000 2.2100 1.2800 2.2100
                 1.2800 1.7200 1.6200 1.7200 1.6200 1.1100 1.5600 1.1100 1.5600 0.6400 1.3200 0.6400
                 1.3200 0.4000 1.4400 0.4000 1.4400 0.5200 1.6800 0.5200 1.6800 0.9900 2.4400 0.9900 ;
        POLYGON  1.5000 1.6000 1.3800 1.6000 1.3800 1.3500 1.3200 1.3500 1.3200 1.0000 1.1200 1.0000
                 1.1200 0.8800 0.2400 0.8800 0.2400 1.8400 0.3200 1.8400 0.3200 2.0800 0.2000 2.0800
                 0.2000 1.9600 0.1200 1.9600 0.1200 0.6400 0.2000 0.6400 0.2000 0.5000 0.3200 0.5000
                 0.3200 0.7600 1.4400 0.7600 1.4400 1.2300 1.5000 1.2300 ;
    END
END CLKMX2X4

MACRO CLKMX2X3
    CLASS CORE ;
    FOREIGN CLKMX2X3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 1.3000 1.5050 1.4200 ;
        RECT  0.4650 1.5200 1.3850 1.6400 ;
        RECT  1.2650 1.3000 1.3850 1.6400 ;
        RECT  0.4650 1.3150 0.5850 1.6400 ;
        RECT  0.3600 1.1950 0.5650 1.4350 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2100 1.1450 1.4000 ;
        RECT  0.7050 1.2100 1.1450 1.3650 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1450 1.2300 2.5950 1.3800 ;
        RECT  2.1450 1.2000 2.2650 1.4400 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4850 1.3150 3.6050 2.2100 ;
        RECT  2.8250 0.7700 3.6050 0.8900 ;
        RECT  3.4850 0.5900 3.6050 0.8900 ;
        RECT  2.8250 1.3150 3.6050 1.4350 ;
        RECT  2.8250 1.1750 3.1200 1.4350 ;
        RECT  2.6450 1.5000 2.9450 1.6200 ;
        RECT  2.8250 0.6500 2.9450 1.6200 ;
        RECT  2.5850 0.6500 2.9450 0.7700 ;
        RECT  2.6450 1.5000 2.7650 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.0650 -0.1800 3.1850 0.6400 ;
        RECT  2.2250 -0.1800 2.3450 0.6400 ;
        RECT  0.6050 -0.1800 0.7250 0.8150 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.0650 1.5600 3.1850 2.7900 ;
        RECT  2.2250 1.5600 2.3450 2.7900 ;
        RECT  0.7650 1.7600 1.0050 2.1500 ;
        RECT  0.7650 1.7600 0.8850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.6850 1.0900 2.4450 1.0900 2.4450 1.0800 2.0250 1.0800 2.0250 1.6800 1.7050 1.6800
                 1.7050 2.2100 1.5850 2.2100 1.5850 1.5600 1.9050 1.5600 1.9050 1.0800 1.8650 1.0800
                 1.8650 0.7700 1.1850 0.7700 1.1850 0.6500 1.9850 0.6500 1.9850 0.9600 2.6850 0.9600 ;
        POLYGON  1.7850 1.4400 1.6650 1.4400 1.6650 1.3200 1.6250 1.3200 1.6250 1.0900 1.0450 1.0900
                 1.0450 1.0550 0.2400 1.0550 0.2400 1.5550 0.3450 1.5550 0.3450 1.8000 0.2250 1.8000
                 0.2250 1.6750 0.1200 1.6750 0.1200 0.8150 0.1850 0.8150 0.1850 0.5750 0.3050 0.5750
                 0.3050 0.9350 1.7450 0.9350 1.7450 1.2000 1.7850 1.2000 ;
    END
END CLKMX2X3

MACRO CLKMX2X2
    CLASS CORE ;
    FOREIGN CLKMX2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.6050 1.1850 1.7250 ;
        RECT  1.0650 1.3100 1.1850 1.7250 ;
        RECT  0.3600 1.4650 0.5100 1.7250 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6450 1.2800 0.8850 1.4850 ;
        RECT  0.6500 1.0900 0.8000 1.4850 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9050 1.2400 2.3050 1.3800 ;
        RECT  2.0450 1.2300 2.3050 1.3800 ;
        RECT  1.9050 1.2400 2.0250 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.1750 2.8300 1.4350 ;
        RECT  2.4250 1.1750 2.8300 1.2950 ;
        RECT  2.4250 0.5900 2.5450 1.6200 ;
        RECT  2.4050 1.5000 2.5250 2.2100 ;
        RECT  2.3450 0.4700 2.4650 0.7100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.7650 -0.1800 2.8850 0.6500 ;
        RECT  1.9250 -0.1800 2.0450 0.7100 ;
        RECT  0.6250 -0.1800 0.7450 0.7100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.8250 1.5600 2.9450 2.7900 ;
        RECT  1.9850 1.8500 2.1050 2.7900 ;
        RECT  0.7050 1.9700 0.8250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3050 1.1000 2.0650 1.1000 2.0650 0.9500 1.7850 0.9500 1.7850 2.0100 1.5250 2.0100
                 1.5250 2.0300 1.2850 2.0300 1.2850 1.9100 1.4050 1.9100 1.4050 1.8900 1.6650 1.8900
                 1.6650 0.9500 1.4250 0.9500 1.4250 0.7300 1.2650 0.7300 1.2650 0.4700 1.3850 0.4700
                 1.3850 0.6100 1.5450 0.6100 1.5450 0.8300 2.3050 0.8300 ;
        POLYGON  1.5450 1.7700 1.4250 1.7700 1.4250 1.1900 1.0650 1.1900 1.0650 0.9700 0.2400 0.9700
                 0.2400 1.8450 0.4050 1.8450 0.4050 2.0900 0.2850 2.0900 0.2850 1.9650 0.1200 1.9650
                 0.1200 0.7300 0.2050 0.7300 0.2050 0.4700 0.3250 0.4700 0.3250 0.8500 1.3050 0.8500
                 1.3050 1.0700 1.5450 1.0700 ;
    END
END CLKMX2X2

MACRO CLKMX2X12
    CLASS CORE ;
    FOREIGN CLKMX2X12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1940  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 1.4150 1.2700 1.5350 ;
        RECT  0.3900 1.5550 1.1100 1.6750 ;
        RECT  0.9900 1.4150 1.1100 1.6750 ;
        RECT  0.3900 1.1750 0.5100 1.6750 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END S0
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0950 0.8700 1.4350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0860  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9300 1.2150 2.2500 1.4350 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.9300 1.2150 2.0500 1.4550 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.9500 1.3100 6.0700 2.2100 ;
        RECT  5.7700 1.3100 6.0700 1.4300 ;
        RECT  5.7900 0.4050 5.9100 1.1600 ;
        RECT  2.6100 1.1900 5.8900 1.3100 ;
        RECT  4.9500 1.0400 5.8900 1.3100 ;
        RECT  5.1100 1.0400 5.2300 2.2100 ;
        RECT  4.9500 0.4050 5.0700 1.3100 ;
        RECT  4.2700 1.1900 4.3900 2.2100 ;
        RECT  3.2700 1.0400 4.2300 1.3100 ;
        RECT  4.1100 0.4050 4.2300 1.3100 ;
        RECT  3.4300 1.0400 3.5500 2.2100 ;
        RECT  3.2700 0.4050 3.3900 1.3100 ;
        RECT  2.6100 1.1750 2.8300 1.4350 ;
        RECT  2.6100 0.6950 2.7300 1.4800 ;
        RECT  2.5900 1.3600 2.7100 2.2100 ;
        RECT  2.3700 0.4600 2.6100 0.8150 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  6.2100 -0.1800 6.3300 0.9200 ;
        RECT  5.3700 -0.1800 5.4900 0.9200 ;
        RECT  4.5300 -0.1800 4.6500 0.9200 ;
        RECT  3.6900 -0.1800 3.8100 0.9200 ;
        RECT  2.8500 -0.1800 2.9700 0.9200 ;
        RECT  1.9500 0.4600 2.1900 0.8150 ;
        RECT  1.9500 -0.1800 2.0700 0.8150 ;
        RECT  0.6100 -0.1800 0.7300 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  6.3700 1.4300 6.4900 2.7900 ;
        RECT  5.5300 1.4300 5.6500 2.7900 ;
        RECT  4.6900 1.4300 4.8100 2.7900 ;
        RECT  3.8500 1.4300 3.9700 2.7900 ;
        RECT  3.0100 1.4300 3.1300 2.7900 ;
        RECT  2.1700 1.5550 2.2900 2.7900 ;
        RECT  0.5900 1.7950 0.7100 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4900 1.2400 2.3700 1.2400 2.3700 1.0550 1.8100 1.0550 1.8100 1.8400 1.4300 1.8400
                 1.4300 2.2100 1.3100 2.2100 1.3100 1.7200 1.6900 1.7200 1.6900 1.0550 1.4100 1.0550
                 1.4100 0.7350 1.2500 0.7350 1.2500 0.4950 1.3700 0.4950 1.3700 0.6150 1.5300 0.6150
                 1.5300 0.9350 2.4900 0.9350 ;
        POLYGON  1.5700 1.6000 1.4500 1.6000 1.4500 1.2950 1.1700 1.2950 1.1700 1.0000 1.0500 1.0000
                 1.0500 0.9750 0.2400 0.9750 0.2400 1.7950 0.2900 1.7950 0.2900 2.2100 0.1700 2.2100
                 0.1700 1.9150 0.1200 1.9150 0.1200 0.7350 0.1900 0.7350 0.1900 0.5900 0.3100 0.5900
                 0.3100 0.8550 1.2900 0.8550 1.2900 1.1750 1.5700 1.1750 ;
    END
END CLKMX2X12

MACRO CLKINVX8
    CLASS CORE ;
    FOREIGN CLKINVX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.8640  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9050 1.2050 2.2650 1.3250 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1450 0.7400 3.3850 0.8600 ;
        RECT  3.2050 1.4700 3.3250 2.2100 ;
        RECT  0.7450 0.7900 3.2650 0.9100 ;
        RECT  0.6850 1.5000 3.3250 1.6200 ;
        RECT  2.3850 0.7900 2.5400 1.1450 ;
        RECT  2.3850 0.7900 2.5050 1.6200 ;
        RECT  2.3650 1.4700 2.4850 2.2100 ;
        RECT  2.3650 0.6700 2.4850 0.9100 ;
        RECT  1.4650 0.7400 1.7050 0.9100 ;
        RECT  1.5250 1.4650 1.6450 2.2100 ;
        RECT  0.6250 0.7400 0.8650 0.8600 ;
        RECT  0.6850 1.5000 0.8050 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.7850 -0.1800 2.9050 0.6700 ;
        RECT  1.9450 -0.1800 2.0650 0.6700 ;
        RECT  1.1050 -0.1800 1.2250 0.6700 ;
        RECT  0.2650 -0.1800 0.3850 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.7850 1.7400 2.9050 2.7900 ;
        RECT  1.9450 1.7400 2.0650 2.7900 ;
        RECT  1.1050 1.7400 1.2250 2.7900 ;
        RECT  0.2650 1.4650 0.3850 2.7900 ;
        END
    END VDD
END CLKINVX8

MACRO CLKINVX6
    CLASS CORE ;
    FOREIGN CLKINVX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8400 1.1500 1.4000 1.2700 ;
        RECT  0.8850 1.1500 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3200 1.4300 2.4400 2.2100 ;
        RECT  0.5800 0.9100 2.4400 1.0300 ;
        RECT  2.3200 0.4000 2.4400 1.0300 ;
        RECT  0.6400 1.5000 2.4400 1.6200 ;
        RECT  1.5200 1.1750 1.6700 1.6200 ;
        RECT  1.5200 0.9100 1.6400 1.6200 ;
        RECT  1.4800 1.4300 1.6000 2.2100 ;
        RECT  1.4800 0.4000 1.6000 1.0300 ;
        RECT  0.6400 1.4300 0.7600 2.2100 ;
        RECT  0.5800 0.4000 0.7000 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.9000 -0.1800 2.0200 0.7900 ;
        RECT  1.0600 -0.1800 1.1800 0.7900 ;
        RECT  0.1600 -0.1800 0.2800 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.9000 1.7400 2.0200 2.7900 ;
        RECT  1.0600 1.7400 1.1800 2.7900 ;
        RECT  0.2200 1.4300 0.3400 2.7900 ;
        END
    END VDD
END CLKINVX6

MACRO CLKINVX4
    CLASS CORE ;
    FOREIGN CLKINVX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8000 1.2600 1.4000 1.3800 ;
        RECT  0.8850 1.2300 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.5200 0.8500 1.6400 1.7250 ;
        RECT  1.5000 1.5000 1.6200 2.2100 ;
        RECT  0.6600 0.8500 1.6400 0.9700 ;
        RECT  1.5000 0.6800 1.6200 0.9700 ;
        RECT  0.6600 1.5000 1.6700 1.6200 ;
        RECT  0.6600 1.5000 0.7800 2.2100 ;
        RECT  0.6600 0.6800 0.7800 0.9700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.9200 -0.1800 2.0400 0.7300 ;
        RECT  1.0800 -0.1800 1.2000 0.7300 ;
        RECT  0.2400 -0.1800 0.3600 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.9200 1.5600 2.0400 2.7900 ;
        RECT  1.0800 1.7400 1.2000 2.7900 ;
        RECT  0.2400 1.5600 0.3600 2.7900 ;
        END
    END VDD
END CLKINVX4

MACRO CLKINVX3
    CLASS CORE ;
    FOREIGN CLKINVX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3240  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.7900 0.4150 1.2450 ;
        RECT  0.2950 0.7600 0.4150 1.2450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.1250 1.5150 2.0150 ;
        RECT  0.6500 0.7600 1.5150 0.8800 ;
        RECT  1.3950 0.5900 1.5150 0.8800 ;
        RECT  0.6500 1.1250 1.5150 1.2450 ;
        RECT  0.6500 0.7600 0.8000 1.2450 ;
        RECT  0.6500 0.7100 0.7700 1.4850 ;
        RECT  0.5550 1.3650 0.6750 2.0150 ;
        RECT  0.5550 0.5900 0.6750 0.8300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.3650 1.0950 2.7900 ;
        RECT  0.1350 1.3650 0.2550 2.7900 ;
        END
    END VDD
END CLKINVX3

MACRO CLKINVX20
    CLASS CORE ;
    FOREIGN CLKINVX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.1600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 1.1650 6.3650 1.2850 ;
        RECT  0.8850 1.1650 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.6132  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2850 1.4500 7.4050 2.2100 ;
        RECT  0.5550 0.9250 7.4050 1.0450 ;
        RECT  7.2850 0.4000 7.4050 1.0450 ;
        RECT  0.5650 1.5000 7.4050 1.6200 ;
        RECT  6.7400 1.1750 6.8900 1.6200 ;
        RECT  6.4850 1.3150 6.8900 1.6200 ;
        RECT  6.4850 0.9250 6.6050 1.6200 ;
        RECT  6.4450 1.4450 6.5650 2.2100 ;
        RECT  6.4450 0.4000 6.5650 1.0450 ;
        RECT  5.6050 1.4450 5.7250 2.2100 ;
        RECT  5.6050 0.4000 5.7250 1.0450 ;
        RECT  4.7650 1.4450 4.8850 2.2100 ;
        RECT  4.7650 0.4000 4.8850 1.0450 ;
        RECT  3.9250 1.4450 4.0450 2.2100 ;
        RECT  3.9250 0.4000 4.0450 1.0450 ;
        RECT  3.0850 1.4450 3.2050 2.2100 ;
        RECT  3.0850 0.4000 3.2050 1.0450 ;
        RECT  2.2450 1.4450 2.3650 2.2100 ;
        RECT  2.2450 0.4000 2.3650 1.0450 ;
        RECT  1.4050 1.4450 1.5250 2.2100 ;
        RECT  1.3950 0.4000 1.5150 1.0450 ;
        RECT  0.5650 1.4450 0.6850 2.2100 ;
        RECT  0.5550 0.4000 0.6750 1.0450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.8650 -0.1800 6.9850 0.8050 ;
        RECT  6.0250 -0.1800 6.1450 0.8050 ;
        RECT  5.1850 -0.1800 5.3050 0.8050 ;
        RECT  4.3450 -0.1800 4.4650 0.8050 ;
        RECT  3.5050 -0.1800 3.6250 0.8050 ;
        RECT  2.6650 -0.1800 2.7850 0.8050 ;
        RECT  1.8250 -0.1800 1.9450 0.8050 ;
        RECT  0.9750 -0.1800 1.0950 0.8050 ;
        RECT  0.1350 -0.1800 0.2550 0.9100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.8650 1.7400 6.9850 2.7900 ;
        RECT  6.0250 1.7400 6.1450 2.7900 ;
        RECT  5.1850 1.7400 5.3050 2.7900 ;
        RECT  4.3450 1.7400 4.4650 2.7900 ;
        RECT  3.5050 1.7400 3.6250 2.7900 ;
        RECT  2.6650 1.7400 2.7850 2.7900 ;
        RECT  1.8250 1.7400 1.9450 2.7900 ;
        RECT  0.9850 1.7400 1.1050 2.7900 ;
        RECT  0.1450 1.4450 0.2650 2.7900 ;
        END
    END VDD
END CLKINVX20

MACRO CLKINVX2
    CLASS CORE ;
    FOREIGN CLKINVX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.4500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3700 1.0000 0.4900 1.2400 ;
        RECT  0.0700 1.0250 0.4900 1.1450 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        RECT  0.6500 0.6800 0.7700 2.0100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.4500 0.1800 ;
        RECT  1.0700 -0.1800 1.1900 0.7300 ;
        RECT  0.2300 -0.1800 0.3500 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.4500 2.7900 ;
        RECT  1.0700 1.3600 1.1900 2.7900 ;
        RECT  0.2300 1.3600 0.3500 2.7900 ;
        END
    END VDD
END CLKINVX2

MACRO CLKINVX16
    CLASS CORE ;
    FOREIGN CLKINVX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.7280  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7750 1.2050 5.4950 1.3250 ;
        RECT  0.8850 1.2050 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5000 5.7350 1.6200 ;
        RECT  5.6150 0.7900 5.7350 1.6200 ;
        RECT  5.5800 1.4650 5.7300 1.7250 ;
        RECT  5.5950 1.4650 5.7150 2.2100 ;
        RECT  0.6150 0.7900 5.7350 0.9100 ;
        RECT  5.5950 0.6700 5.7150 0.9100 ;
        RECT  4.6950 0.7400 4.9350 0.9100 ;
        RECT  4.7550 1.4700 4.8750 2.2100 ;
        RECT  3.8550 0.7400 4.0950 0.9100 ;
        RECT  3.9150 1.4700 4.0350 2.2100 ;
        RECT  3.0150 0.7400 3.2550 0.9100 ;
        RECT  3.0750 1.4650 3.1950 2.2100 ;
        RECT  2.1750 0.7400 2.4150 0.9100 ;
        RECT  2.2350 1.4650 2.3550 2.2100 ;
        RECT  1.3350 0.7400 1.5750 0.9100 ;
        RECT  1.3950 1.4650 1.5150 2.2100 ;
        RECT  0.4950 0.7400 0.7350 0.8600 ;
        RECT  0.5550 1.4650 0.6750 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  6.0150 -0.1800 6.1350 0.6700 ;
        RECT  5.1750 -0.1800 5.2950 0.6700 ;
        RECT  4.3350 -0.1800 4.4550 0.6700 ;
        RECT  3.4950 -0.1800 3.6150 0.6700 ;
        RECT  2.6550 -0.1800 2.7750 0.6700 ;
        RECT  1.8150 -0.1800 1.9350 0.6700 ;
        RECT  0.9750 -0.1800 1.0950 0.6650 ;
        RECT  0.1350 -0.1800 0.2550 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  6.0150 1.4700 6.1350 2.7900 ;
        RECT  5.1750 1.7400 5.2950 2.7900 ;
        RECT  4.3350 1.7400 4.4550 2.7900 ;
        RECT  3.4950 1.7400 3.6150 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.4650 0.2550 2.7900 ;
        END
    END VDD
END CLKINVX16

MACRO CLKINVX12
    CLASS CORE ;
    FOREIGN CLKINVX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.2960  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 1.1500 3.8350 1.2700 ;
        RECT  0.8850 1.1500 1.1450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.5000 4.0750 1.6200 ;
        RECT  3.9550 0.9100 4.0750 1.6200 ;
        RECT  3.9150 1.4300 4.0350 2.2100 ;
        RECT  0.5550 0.9100 4.0750 1.0300 ;
        RECT  3.9150 0.4000 4.0350 1.0300 ;
        RECT  3.8400 1.4650 4.0350 1.7250 ;
        RECT  3.0750 1.4300 3.1950 2.2100 ;
        RECT  3.0750 0.4000 3.1950 1.0300 ;
        RECT  2.2350 1.4300 2.3550 2.2100 ;
        RECT  2.2350 0.4000 2.3550 1.0300 ;
        RECT  1.3950 1.4300 1.5150 2.2100 ;
        RECT  1.3950 0.4000 1.5150 1.0300 ;
        RECT  0.5550 1.4300 0.6750 2.2100 ;
        RECT  0.5550 0.4000 0.6750 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  4.3350 -0.1800 4.4550 0.9150 ;
        RECT  3.4950 -0.1800 3.6150 0.7900 ;
        RECT  2.6550 -0.1800 2.7750 0.7900 ;
        RECT  1.8150 -0.1800 1.9350 0.7900 ;
        RECT  0.9750 -0.1800 1.0950 0.7900 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  4.3350 1.4300 4.4550 2.7900 ;
        RECT  3.4950 1.7400 3.6150 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.4300 0.2550 2.7900 ;
        END
    END VDD
END CLKINVX12

MACRO CLKINVX1
    CLASS CORE ;
    FOREIGN CLKINVX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 0.8700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 0.7950 0.2400 1.2200 ;
        RECT  0.0700 0.7950 0.2400 1.2000 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 0.6250 0.6750 1.9900 ;
        RECT  0.3600 0.8850 0.6750 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 0.8700 0.1800 ;
        RECT  0.1350 -0.1800 0.2550 0.6750 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 0.8700 2.7900 ;
        RECT  0.1350 1.3400 0.2550 2.7900 ;
        END
    END VDD
END CLKINVX1

MACRO CLKBUFX8
    CLASS CORE ;
    FOREIGN CLKBUFX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8700 0.8250 3.9900 1.3050 ;
        RECT  3.8400 0.8250 3.9900 1.2800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6900 0.7150 2.9300 0.8350 ;
        RECT  2.7500 1.2950 2.8700 2.2100 ;
        RECT  0.2300 0.7600 2.8100 0.8800 ;
        RECT  2.5700 1.2950 2.8700 1.4150 ;
        RECT  0.2300 1.2700 2.6900 1.3900 ;
        RECT  1.8500 0.7100 2.0900 0.8800 ;
        RECT  1.9100 1.2700 2.0300 2.2100 ;
        RECT  1.0100 0.7100 1.2500 0.8800 ;
        RECT  1.0700 1.2700 1.1900 2.2100 ;
        RECT  0.3600 0.7600 0.5100 1.1450 ;
        RECT  0.3600 0.7600 0.4800 1.3900 ;
        RECT  0.2300 1.2700 0.3500 2.2100 ;
        RECT  0.2300 0.6400 0.3500 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  4.0100 -0.1800 4.1300 0.7050 ;
        RECT  3.1700 -0.1800 3.2900 0.7050 ;
        RECT  2.3300 -0.1800 2.4500 0.6400 ;
        RECT  1.4900 -0.1800 1.6100 0.6400 ;
        RECT  0.6500 -0.1800 0.7700 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  4.0100 1.4650 4.1300 2.7900 ;
        RECT  3.1700 1.4650 3.2900 2.7900 ;
        RECT  2.3300 1.5100 2.4500 2.7900 ;
        RECT  1.4900 1.5100 1.6100 2.7900 ;
        RECT  0.6500 1.5100 0.7700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.7100 2.1150 3.5900 2.1150 3.5900 1.1500 3.1900 1.1500 3.1900 1.1750 2.9500 1.1750
                 2.9500 1.1500 0.8700 1.1500 0.8700 1.0300 3.5900 1.0300 3.5900 0.6550 3.7100 0.6550 ;
    END
END CLKBUFX8

MACRO CLKBUFX6
    CLASS CORE ;
    FOREIGN CLKBUFX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8900 1.3900 2.0100 2.2100 ;
        RECT  0.1500 0.9100 2.0100 1.0300 ;
        RECT  1.8900 0.4000 2.0100 1.0300 ;
        RECT  0.2100 1.3900 2.0100 1.5100 ;
        RECT  1.0500 1.3900 1.1700 2.2100 ;
        RECT  0.9900 0.4000 1.1100 1.0300 ;
        RECT  0.3600 1.1750 0.5100 1.5100 ;
        RECT  0.3600 0.9100 0.4800 1.5100 ;
        RECT  0.2100 1.3900 0.3300 2.2100 ;
        RECT  0.1500 0.4000 0.2700 1.0300 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.8250 3.1200 1.2850 ;
        RECT  2.9700 0.8250 3.0900 1.3100 ;
        END
    END A
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  3.1500 1.4300 3.2700 2.7900 ;
        RECT  2.3100 1.4300 2.4300 2.7900 ;
        RECT  1.4700 1.6300 1.5900 2.7900 ;
        RECT  0.6300 1.6300 0.7500 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  3.1500 -0.1800 3.2700 0.7050 ;
        RECT  2.3100 -0.1800 2.4300 0.8950 ;
        RECT  1.4100 -0.1800 1.5300 0.7900 ;
        RECT  0.5700 -0.1800 0.6900 0.7900 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  2.8500 2.0800 2.7300 2.0800 2.7300 1.2700 0.7700 1.2700 0.7700 1.1500 2.7300 1.1500
                 2.7300 0.6550 2.8500 0.6550 ;
    END
END CLKBUFX6

MACRO CLKBUFX4
    CLASS CORE ;
    FOREIGN CLKBUFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9550 1.2400 2.0750 1.4800 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.8400 1.3600 2.0750 1.4800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3350 0.7100 1.5750 0.8300 ;
        RECT  1.3950 1.3200 1.5150 2.2100 ;
        RECT  0.5150 0.7600 1.4550 0.8800 ;
        RECT  0.5150 1.3200 1.5150 1.4400 ;
        RECT  0.5550 1.3200 0.8000 1.7250 ;
        RECT  0.5550 1.3200 0.6750 2.2100 ;
        RECT  0.5550 0.6400 0.6750 0.8800 ;
        RECT  0.5150 0.7600 0.6350 1.4400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8150 -0.1800 1.9350 0.7000 ;
        RECT  0.9150 0.5200 1.1550 0.6400 ;
        RECT  0.9150 -0.1800 1.0350 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8150 1.8450 1.9350 2.7900 ;
        RECT  0.9750 1.5600 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3550 2.2100 2.2350 2.2100 2.2350 1.1200 1.4150 1.1200 1.4150 1.1700 1.1750 1.1700
                 1.1750 1.1200 0.9950 1.1200 0.9950 1.1700 0.7550 1.1700 0.7550 1.0500 0.8750 1.0500
                 0.8750 1.0000 2.2350 1.0000 2.2350 0.6500 2.3550 0.6500 ;
    END
END CLKBUFX4

MACRO CLKBUFX3
    CLASS CORE ;
    FOREIGN CLKBUFX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.0000 1.6700 1.5000 ;
        RECT  1.5200 1.0000 1.6700 1.4700 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9750 1.3200 1.0950 2.2100 ;
        RECT  0.9750 0.4000 1.0950 0.6400 ;
        RECT  0.1350 0.7600 1.0900 0.8800 ;
        RECT  0.1350 1.3200 1.0950 1.4400 ;
        RECT  0.9700 0.5200 1.0900 0.8800 ;
        RECT  0.3600 1.1750 0.5100 1.4400 ;
        RECT  0.3600 0.7600 0.4800 1.4400 ;
        RECT  0.1350 1.3200 0.2550 2.2100 ;
        RECT  0.1350 0.5900 0.2550 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.3950 1.6200 1.5150 2.7900 ;
        RECT  0.5550 1.5600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 2.2100 1.8150 2.2100 1.8150 0.8800 1.3300 0.8800 1.3300 1.1700 1.2100 1.1700
                 1.2100 0.7600 1.8150 0.7600 1.8150 0.5900 1.9350 0.5900 ;
    END
END CLKBUFX3

MACRO CLKBUFX20
    CLASS CORE ;
    FOREIGN CLKBUFX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.5400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0200 1.2600 8.6200 1.3800 ;
        RECT  8.1350 1.2300 8.3950 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.6387  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9600 1.4250 7.0800 2.2100 ;
        RECT  0.3600 0.9450 7.0800 1.0650 ;
        RECT  6.9600 0.4000 7.0800 1.0650 ;
        RECT  0.2400 1.4250 7.0800 1.5450 ;
        RECT  6.1200 1.4250 6.2400 2.2100 ;
        RECT  6.1200 0.4000 6.2400 1.0650 ;
        RECT  5.2800 1.4250 5.4000 2.2100 ;
        RECT  5.2200 0.4000 5.3400 1.0650 ;
        RECT  4.4400 1.4250 4.5600 2.2100 ;
        RECT  4.3800 0.4000 4.5000 1.0650 ;
        RECT  3.6000 1.4250 3.7200 2.2100 ;
        RECT  3.5400 0.4000 3.6600 1.0650 ;
        RECT  2.7600 1.4250 2.8800 2.2100 ;
        RECT  2.7000 0.4000 2.8200 1.0650 ;
        RECT  1.9200 1.4250 2.0400 2.2100 ;
        RECT  1.8600 0.4000 1.9800 1.0650 ;
        RECT  1.0800 1.4250 1.2000 2.2100 ;
        RECT  1.0200 0.4000 1.1400 1.0650 ;
        RECT  0.3600 0.9450 0.5100 1.5450 ;
        RECT  0.3600 0.7850 0.4800 1.5450 ;
        RECT  0.2400 1.4250 0.3600 2.2100 ;
        RECT  0.1800 0.7850 0.4800 0.9050 ;
        RECT  0.1800 0.4000 0.3000 0.9050 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.0600 -0.1800 9.1800 0.7200 ;
        RECT  8.2200 -0.1800 8.3400 0.7200 ;
        RECT  7.3800 -0.1800 7.5000 0.9100 ;
        RECT  6.5400 -0.1800 6.6600 0.8250 ;
        RECT  5.6400 -0.1800 5.7600 0.8250 ;
        RECT  4.8000 -0.1800 4.9200 0.8250 ;
        RECT  3.9600 -0.1800 4.0800 0.8250 ;
        RECT  3.1200 -0.1800 3.2400 0.8250 ;
        RECT  2.2800 -0.1800 2.4000 0.8250 ;
        RECT  1.4400 -0.1800 1.5600 0.8250 ;
        RECT  0.6000 -0.1800 0.7200 0.8250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  9.0600 1.7400 9.1800 2.7900 ;
        RECT  8.2200 1.7400 8.3400 2.7900 ;
        RECT  7.3800 1.5600 7.5000 2.7900 ;
        RECT  6.5400 1.6650 6.6600 2.7900 ;
        RECT  5.7000 1.6650 5.8200 2.7900 ;
        RECT  4.8600 1.6650 4.9800 2.7900 ;
        RECT  4.0200 1.6650 4.1400 2.7900 ;
        RECT  3.1800 1.6650 3.3000 2.7900 ;
        RECT  2.3400 1.6650 2.4600 2.7900 ;
        RECT  1.5000 1.6650 1.6200 2.7900 ;
        RECT  0.6600 1.6650 0.7800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.6000 0.9600 7.9000 0.9600 7.9000 1.5000 9.6000 1.5000 9.6000 2.2100 9.4800 2.2100
                 9.4800 1.6200 8.7600 1.6200 8.7600 2.2100 8.6400 2.2100 8.6400 1.6200 7.9200 1.6200
                 7.9200 2.2100 7.8000 2.2100 7.8000 1.6200 7.7800 1.6200 7.7800 1.3050 0.8200 1.3050
                 0.8200 1.1850 7.7800 1.1850 7.7800 0.8400 7.8000 0.8400 7.8000 0.6700 7.9200 0.6700
                 7.9200 0.8400 8.6400 0.8400 8.6400 0.6700 8.7600 0.6700 8.7600 0.8400 9.4800 0.8400
                 9.4800 0.6700 9.6000 0.6700 ;
    END
END CLKBUFX20

MACRO CLKBUFX2
    CLASS CORE ;
    FOREIGN CLKBUFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2250 1.2750 1.3800 ;
        RECT  1.1550 1.1300 1.2750 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.2250 0.6750 2.1200 ;
        RECT  0.5550 0.6050 0.6750 0.8450 ;
        RECT  0.5150 0.7250 0.6350 1.3450 ;
        RECT  0.3600 0.8850 0.6350 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.7700 ;
        RECT  0.1350 -0.1800 0.2550 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.5000 1.0950 2.7900 ;
        RECT  0.1350 1.4700 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5150 1.7400 1.3950 1.7400 1.3950 1.0100 1.0350 1.0100 1.0350 1.1050 0.7550 1.1050
                 0.7550 0.9850 0.9150 0.9850 0.9150 0.8900 1.3950 0.8900 1.3950 0.5300 1.5150 0.5300 ;
    END
END CLKBUFX2

MACRO CLKBUFX16
    CLASS CORE ;
    FOREIGN CLKBUFX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6850 1.2600 7.2850 1.3800 ;
        RECT  6.6850 1.2300 6.9450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5650 0.7150 5.8050 0.8350 ;
        RECT  5.6250 1.2950 5.7450 2.2100 ;
        RECT  0.5450 0.7650 5.6850 0.8850 ;
        RECT  0.5450 1.2950 5.7450 1.4150 ;
        RECT  4.7250 0.7150 4.9650 0.8850 ;
        RECT  4.7850 1.2950 4.9050 2.2100 ;
        RECT  3.8850 0.7150 4.1250 0.8850 ;
        RECT  3.9450 1.2950 4.0650 2.2100 ;
        RECT  3.0450 0.7150 3.2850 0.8850 ;
        RECT  3.1050 1.2950 3.2250 2.2100 ;
        RECT  2.2050 0.7150 2.4450 0.8850 ;
        RECT  2.2650 1.2950 2.3850 2.2100 ;
        RECT  1.3650 0.7150 1.6050 0.8850 ;
        RECT  1.4250 1.2950 1.5450 2.2100 ;
        RECT  0.5850 1.2950 0.8000 1.7250 ;
        RECT  0.5850 1.2950 0.7050 2.2100 ;
        RECT  0.5850 0.6450 0.7050 0.8850 ;
        RECT  0.5450 0.7650 0.6650 1.4150 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.7250 -0.1800 7.8450 0.7050 ;
        RECT  6.8850 -0.1800 7.0050 0.7050 ;
        RECT  6.0450 -0.1800 6.1650 0.7050 ;
        RECT  5.2050 -0.1800 5.3250 0.6450 ;
        RECT  4.3650 -0.1800 4.4850 0.6450 ;
        RECT  3.5250 -0.1800 3.6450 0.6450 ;
        RECT  2.6850 -0.1800 2.8050 0.6450 ;
        RECT  1.8450 -0.1800 1.9650 0.6450 ;
        RECT  1.0050 -0.1800 1.1250 0.6400 ;
        RECT  0.1650 -0.1800 0.2850 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.7250 1.5600 7.8450 2.7900 ;
        RECT  6.8850 1.7400 7.0050 2.7900 ;
        RECT  6.0450 1.5600 6.1650 2.7900 ;
        RECT  5.2050 1.5350 5.3250 2.7900 ;
        RECT  4.3650 1.5350 4.4850 2.7900 ;
        RECT  3.5250 1.5350 3.6450 2.7900 ;
        RECT  2.6850 1.5350 2.8050 2.7900 ;
        RECT  1.8450 1.5350 1.9650 2.7900 ;
        RECT  1.0050 1.5350 1.1250 2.7900 ;
        RECT  0.1650 1.4650 0.2850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.4250 0.9450 6.5650 0.9450 6.5650 1.5000 7.4250 1.5000 7.4250 2.2100 7.3050 2.2100
                 7.3050 1.6200 6.5850 1.6200 6.5850 2.2100 6.4650 2.2100 6.4650 1.6200 6.4450 1.6200
                 6.4450 1.1750 0.7850 1.1750 0.7850 1.0550 6.4450 1.0550 6.4450 0.8250 6.4650 0.8250
                 6.4650 0.6550 6.5850 0.6550 6.5850 0.8250 7.3050 0.8250 7.3050 0.6550 7.4250 0.6550 ;
    END
END CLKBUFX16

MACRO CLKBUFX12
    CLASS CORE ;
    FOREIGN CLKBUFX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3240  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4500 1.3000 4.7750 1.4200 ;
        RECT  4.4200 1.4650 4.5700 1.7250 ;
        RECT  4.4500 1.3000 4.5700 1.7250 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9150 1.3200 4.0350 2.2100 ;
        RECT  0.5150 0.8200 4.0350 0.9400 ;
        RECT  3.9150 0.4000 4.0350 0.9400 ;
        RECT  0.5150 1.3200 4.0350 1.4400 ;
        RECT  3.0750 1.3200 3.1950 2.2100 ;
        RECT  3.0750 0.4000 3.1950 0.9400 ;
        RECT  2.2350 1.3200 2.3550 2.2100 ;
        RECT  2.2350 0.4000 2.3550 0.9400 ;
        RECT  1.3950 1.3200 1.5150 2.2100 ;
        RECT  1.3950 0.4000 1.5150 0.9400 ;
        RECT  0.5550 1.3200 0.8000 1.7250 ;
        RECT  0.5550 1.3200 0.6750 2.2100 ;
        RECT  0.5550 0.4000 0.6750 0.9400 ;
        RECT  0.5150 0.8000 0.6350 1.4400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.1750 -0.1800 5.2950 0.7250 ;
        RECT  4.3350 -0.1800 4.4550 0.9150 ;
        RECT  3.4950 -0.1800 3.6150 0.7000 ;
        RECT  2.6550 -0.1800 2.7750 0.7000 ;
        RECT  1.8150 -0.1800 1.9350 0.7000 ;
        RECT  0.9750 -0.1800 1.0950 0.7000 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1750 1.5600 5.2950 2.7900 ;
        RECT  4.3350 1.8450 4.4550 2.7900 ;
        RECT  3.4950 1.5600 3.6150 2.7900 ;
        RECT  2.6550 1.5600 2.7750 2.7900 ;
        RECT  1.8150 1.5600 1.9350 2.7900 ;
        RECT  0.9750 1.5600 1.0950 2.7900 ;
        RECT  0.1350 1.4300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7150 0.9650 5.0150 0.9650 5.0150 1.3200 5.7150 1.3200 5.7150 2.2100 5.5950 2.2100
                 5.5950 1.4400 5.0150 1.4400 5.0150 1.6600 4.8750 1.6600 4.8750 2.2100 4.7550 2.2100
                 4.7550 1.5400 4.8950 1.5400 4.8950 1.1800 3.9350 1.1800 3.9350 1.1950 3.6950 1.1950
                 3.6950 1.1800 3.0950 1.1800 3.0950 1.1950 2.8550 1.1950 2.8550 1.1800 2.6750 1.1800
                 2.6750 1.1950 2.4350 1.1950 2.4350 1.1800 1.8350 1.1800 1.8350 1.1950 1.5950 1.1950
                 1.5950 1.1800 0.9950 1.1800 0.9950 1.2000 0.7550 1.2000 0.7550 1.0800 0.8750 1.0800
                 0.8750 1.0600 4.7550 1.0600 4.7550 0.6750 4.8750 0.6750 4.8750 0.8450 5.5950 0.8450
                 5.5950 0.6750 5.7150 0.6750 ;
    END
END CLKBUFX12

MACRO CLKAND2X8
    CLASS CORE ;
    FOREIGN CLKAND2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.6700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3020  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1150 0.9650 3.2350 1.2350 ;
        RECT  0.5950 0.9650 3.2350 1.0850 ;
        RECT  1.5950 0.9650 1.8350 1.1150 ;
        RECT  0.4150 1.0150 0.8550 1.1350 ;
        RECT  0.5950 0.9400 0.8550 1.1350 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3020  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.2050 2.5350 1.3250 ;
        RECT  2.0450 1.2050 2.3050 1.3800 ;
        RECT  1.2950 1.2350 2.3050 1.3550 ;
        RECT  1.1750 1.2050 1.4150 1.3250 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4150 1.2950 6.5350 2.2100 ;
        RECT  6.2750 0.7150 6.5150 0.8350 ;
        RECT  3.8950 1.2950 6.5350 1.4150 ;
        RECT  3.8150 0.7650 6.3950 0.8850 ;
        RECT  5.5800 1.1750 5.7300 1.4350 ;
        RECT  5.5800 0.7150 5.7000 1.4350 ;
        RECT  5.5750 1.2950 5.6950 2.2100 ;
        RECT  5.4350 0.7150 5.7000 0.8850 ;
        RECT  4.7350 1.2950 4.8550 2.2100 ;
        RECT  4.5950 0.7150 4.8350 0.8850 ;
        RECT  3.8950 1.2950 4.0150 2.2100 ;
        RECT  3.6950 0.7150 3.9350 0.8350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.6700 0.1800 ;
        RECT  5.9150 -0.1800 6.0350 0.6450 ;
        RECT  5.0750 -0.1800 5.1950 0.6450 ;
        RECT  4.1750 -0.1800 4.2950 0.6400 ;
        RECT  3.2750 0.4600 3.5150 0.5800 ;
        RECT  3.2750 -0.1800 3.3950 0.5800 ;
        RECT  1.7350 0.4850 1.9750 0.6050 ;
        RECT  1.7350 -0.1800 1.8550 0.6050 ;
        RECT  0.3150 -0.1800 0.4350 0.6650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.6700 2.7900 ;
        RECT  5.9950 1.5350 6.1150 2.7900 ;
        RECT  5.1550 1.5350 5.2750 2.7900 ;
        RECT  4.3150 1.5350 4.4350 2.7900 ;
        RECT  3.4150 2.0700 3.5350 2.7900 ;
        RECT  2.6950 2.0700 2.8150 2.7900 ;
        RECT  1.8550 2.0700 1.9750 2.7900 ;
        RECT  1.0150 2.0700 1.1350 2.7900 ;
        RECT  0.1350 2.0700 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.4600 1.1750 3.4750 1.1750 3.4750 1.6450 0.4750 1.6450 0.4750 1.5250 3.3550 1.5250
                 3.3550 0.8450 1.2150 0.8450 1.2150 0.7950 1.0950 0.7950 1.0950 0.6750 1.3350 0.6750
                 1.3350 0.7250 2.5750 0.7250 2.5750 0.6750 2.8150 0.6750 2.8150 0.7250 3.4750 0.7250
                 3.4750 1.0550 5.4600 1.0550 ;
    END
END CLKAND2X8

MACRO CLKAND2X6
    CLASS CORE ;
    FOREIGN CLKAND2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.8000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3020  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1050 0.9400 3.2250 1.2400 ;
        RECT  0.5950 0.9400 3.2250 1.0600 ;
        RECT  1.5350 0.9400 1.7750 1.1100 ;
        RECT  0.3850 0.9900 0.8550 1.1100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3020  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 1.1800 2.5050 1.3000 ;
        RECT  1.7550 1.2300 2.0150 1.3800 ;
        RECT  1.2950 1.2300 2.0150 1.3500 ;
        RECT  1.1450 1.1800 1.4150 1.3000 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5450 1.3900 5.6650 2.2100 ;
        RECT  3.8650 1.3900 5.6650 1.5100 ;
        RECT  5.4050 0.4000 5.5250 0.9150 ;
        RECT  5.2250 0.7950 5.5250 0.9150 ;
        RECT  3.6650 0.9100 5.3450 1.0300 ;
        RECT  4.7450 1.1750 5.1500 1.5100 ;
        RECT  4.7450 0.7950 4.8650 1.5100 ;
        RECT  4.7050 1.3900 4.8250 2.2100 ;
        RECT  4.5650 0.7950 4.8650 1.0300 ;
        RECT  4.5650 0.4000 4.6850 1.0300 ;
        RECT  3.8650 1.3900 3.9850 2.2100 ;
        RECT  3.6650 0.4000 3.7850 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.8000 0.1800 ;
        RECT  4.9850 -0.1800 5.1050 0.7900 ;
        RECT  4.1450 -0.1800 4.2650 0.7900 ;
        RECT  3.1850 0.4600 3.4250 0.5800 ;
        RECT  3.1850 -0.1800 3.3050 0.5800 ;
        RECT  1.6950 0.4600 1.9350 0.5800 ;
        RECT  1.6950 -0.1800 1.8150 0.5800 ;
        RECT  0.2850 -0.1800 0.4050 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.8000 2.7900 ;
        RECT  5.1250 1.6300 5.2450 2.7900 ;
        RECT  4.2850 1.6300 4.4050 2.7900 ;
        RECT  3.3850 2.0450 3.5050 2.7900 ;
        RECT  2.5450 2.0450 2.6650 2.7900 ;
        RECT  1.8250 2.0450 1.9450 2.7900 ;
        RECT  0.9850 2.0450 1.1050 2.7900 ;
        RECT  0.1350 2.0450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.6250 1.2700 3.4650 1.2700 3.4650 1.6200 0.4450 1.6200 0.4450 1.5000 3.3450 1.5000
                 3.3450 0.8200 1.1750 0.8200 1.1750 0.7700 1.0550 0.7700 1.0550 0.6500 1.2950 0.6500
                 1.2950 0.7000 2.5450 0.7000 2.5450 0.6500 2.7850 0.6500 2.7850 0.7000 3.4650 0.7000
                 3.4650 1.1500 4.6250 1.1500 ;
    END
END CLKAND2X6

MACRO CLKAND2X4
    CLASS CORE ;
    FOREIGN CLKAND2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1510  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 1.0400 1.5900 1.1600 ;
        RECT  0.5950 0.9900 1.3850 1.1100 ;
        RECT  0.5950 0.9400 0.8550 1.1100 ;
        RECT  0.3900 1.0400 0.7150 1.1600 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1510  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8350 1.2550 1.1450 1.4800 ;
        RECT  0.8850 1.2300 1.1450 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0300 1.2900 3.1500 2.1800 ;
        RECT  2.9700 1.1750 3.1200 1.4350 ;
        RECT  2.9700 0.7600 3.0900 1.4350 ;
        RECT  2.1900 1.2900 3.1500 1.4100 ;
        RECT  1.9900 0.8100 3.0900 0.9300 ;
        RECT  2.8300 0.7600 3.0900 0.9300 ;
        RECT  2.8300 0.6400 2.9500 0.9300 ;
        RECT  2.1900 1.2900 2.3100 2.1800 ;
        RECT  1.9900 0.6400 2.1100 0.9300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.2500 -0.1800 3.3700 0.6900 ;
        RECT  2.4100 -0.1800 2.5300 0.6900 ;
        RECT  1.5100 0.5100 1.7500 0.6300 ;
        RECT  1.5100 -0.1800 1.6300 0.6300 ;
        RECT  0.2900 -0.1800 0.4100 0.6900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.4500 1.5300 3.5700 2.7900 ;
        RECT  2.6100 1.5300 2.7300 2.7900 ;
        RECT  1.7100 2.1350 1.8300 2.7900 ;
        RECT  0.8700 2.1350 0.9900 2.7900 ;
        RECT  0.1350 2.1350 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.8500 1.1700 1.8300 1.1700 1.8300 1.7200 0.4500 1.7200 0.4500 1.6000 1.7100 1.6000
                 1.7100 0.8700 0.9900 0.8700 0.9900 0.8200 0.8700 0.8200 0.8700 0.7000 1.1100 0.7000
                 1.1100 0.7500 1.8300 0.7500 1.8300 1.0500 2.8500 1.0500 ;
    END
END CLKAND2X4

MACRO CLKAND2X3
    CLASS CORE ;
    FOREIGN CLKAND2X3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1510  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2650 1.0200 1.6650 1.1400 ;
        RECT  0.5950 0.9700 1.3850 1.0900 ;
        RECT  0.5950 0.9400 0.8550 1.0900 ;
        RECT  0.4350 1.0200 0.7650 1.1400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1510  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2100 1.1450 1.4800 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2250 1.2500 3.3450 2.1400 ;
        RECT  2.3900 1.2500 3.3450 1.3700 ;
        RECT  2.2650 0.7900 3.0450 0.9100 ;
        RECT  2.9250 0.6200 3.0450 0.9100 ;
        RECT  2.3900 0.7900 2.5400 1.3700 ;
        RECT  2.3850 1.2700 2.5100 1.3900 ;
        RECT  2.3850 1.2700 2.5050 2.1400 ;
        RECT  2.0250 0.6800 2.3850 0.8000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.5050 -0.1800 2.6250 0.6700 ;
        RECT  1.6050 0.4900 1.8450 0.6100 ;
        RECT  1.6050 -0.1800 1.7250 0.6100 ;
        RECT  0.3350 -0.1800 0.4550 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  2.8050 1.4900 2.9250 2.7900 ;
        RECT  1.9050 2.0950 2.0250 2.7900 ;
        RECT  1.0350 2.0950 1.1550 2.7900 ;
        RECT  0.1350 1.5750 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2700 1.1500 1.9050 1.1500 1.9050 1.7200 0.4950 1.7200 0.4950 1.6000 1.7850 1.6000
                 1.7850 0.8500 1.0650 0.8500 1.0650 0.8000 0.9450 0.8000 0.9450 0.6800 1.1850 0.6800
                 1.1850 0.7300 1.9050 0.7300 1.9050 1.0300 2.2700 1.0300 ;
    END
END CLKAND2X3

MACRO CLKAND2X2
    CLASS CORE ;
    FOREIGN CLKAND2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0840  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2350 1.2350 0.3550 1.4750 ;
        RECT  0.0700 1.2350 0.3550 1.4350 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0840  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.7750 1.1750 1.0900 1.2950 ;
        RECT  0.7750 1.0550 0.8950 1.2950 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4500 0.8850 1.6700 1.1450 ;
        RECT  1.4500 0.5750 1.5700 1.4450 ;
        RECT  1.3550 1.3250 1.4750 2.0450 ;
        RECT  1.3550 0.4550 1.4750 0.6950 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  1.7750 -0.1800 1.8950 0.6950 ;
        RECT  0.8750 -0.1800 0.9950 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.7750 1.3950 1.8950 2.7900 ;
        RECT  0.9350 1.5550 1.0550 2.7900 ;
        RECT  0.1350 2.1950 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.3300 1.2050 1.2100 1.2050 1.2100 0.9350 0.6350 0.9350 0.6350 1.7950 0.5150 1.7950
                 0.5150 0.8600 0.1750 0.8600 0.1750 0.7400 0.6350 0.7400 0.6350 0.8150 1.3300 0.8150 ;
    END
END CLKAND2X2

MACRO CLKAND2X12
    CLASS CORE ;
    FOREIGN CLKAND2X12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4530  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2550 1.0000 3.3750 1.2400 ;
        RECT  0.6800 1.0000 3.3750 1.1200 ;
        RECT  1.9900 1.0000 2.2300 1.1950 ;
        RECT  0.6500 1.0750 0.8000 1.4350 ;
        RECT  0.4350 1.0750 0.8000 1.1950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4530  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4950 1.2800 4.2550 1.4000 ;
        RECT  1.2700 1.3600 3.7550 1.4800 ;
        RECT  3.4950 1.2300 3.7550 1.4800 ;
        RECT  2.3900 1.2400 2.5100 1.4800 ;
        RECT  1.2700 1.2400 1.3900 1.4800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2500 1.3900 8.3700 2.2100 ;
        RECT  8.1900 1.1750 8.3400 1.5100 ;
        RECT  8.1900 0.7950 8.3100 1.5100 ;
        RECT  4.8900 1.3900 8.3700 1.5100 ;
        RECT  4.6550 0.9100 8.3100 1.0300 ;
        RECT  8.0500 0.7950 8.3100 1.0300 ;
        RECT  8.0500 0.4000 8.1700 1.0300 ;
        RECT  7.4100 1.3900 7.5300 2.2100 ;
        RECT  7.2100 0.4000 7.3300 1.0300 ;
        RECT  6.5700 1.3900 6.6900 2.2100 ;
        RECT  6.3700 0.4000 6.4900 1.0300 ;
        RECT  5.7300 1.3900 5.8500 2.2100 ;
        RECT  5.5300 0.4000 5.6500 1.0300 ;
        RECT  4.8900 1.3900 5.0100 2.2100 ;
        RECT  4.6550 0.4000 4.7750 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.4700 -0.1800 8.5900 0.9150 ;
        RECT  7.6300 -0.1800 7.7500 0.7900 ;
        RECT  6.7900 -0.1800 6.9100 0.7900 ;
        RECT  5.9500 -0.1800 6.0700 0.7900 ;
        RECT  5.0750 -0.1800 5.1950 0.7900 ;
        RECT  4.2350 -0.1800 4.3550 0.6400 ;
        RECT  2.5300 -0.1800 2.6500 0.6400 ;
        RECT  0.9900 -0.1800 1.1100 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.6700 1.4300 8.7900 2.7900 ;
        RECT  7.8300 1.6300 7.9500 2.7900 ;
        RECT  6.9900 1.6300 7.1100 2.7900 ;
        RECT  6.1500 1.6300 6.2700 2.7900 ;
        RECT  5.3100 1.6300 5.4300 2.7900 ;
        RECT  4.4100 2.2300 4.5300 2.7900 ;
        RECT  3.5700 2.2300 3.6900 2.7900 ;
        RECT  2.7300 2.2300 2.8500 2.7900 ;
        RECT  1.8900 2.2300 2.0100 2.7900 ;
        RECT  1.0350 2.2300 1.1550 2.7900 ;
        RECT  0.1350 1.7100 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.0700 1.2700 4.4950 1.2700 4.4950 1.7400 0.4950 1.7400 0.4950 1.6200 4.3750 1.6200
                 4.3750 0.8800 3.7150 0.8800 3.7150 0.9200 3.5950 0.9200 3.5950 0.8800 0.4550 0.8800
                 0.4550 0.9150 0.3350 0.9150 0.3350 0.4000 0.4550 0.4000 0.4550 0.7600 1.7900 0.7600
                 1.7900 0.4000 1.9100 0.4000 1.9100 0.7600 3.5950 0.7600 3.5950 0.4000 3.7150 0.4000
                 3.7150 0.7600 4.4950 0.7600 4.4950 1.1500 8.0700 1.1500 ;
    END
END CLKAND2X12

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8700 0.8250 3.9900 1.3050 ;
        RECT  3.8400 0.8250 3.9900 1.2800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6900 0.7150 2.9300 0.8350 ;
        RECT  2.7500 1.2950 2.8700 2.2100 ;
        RECT  0.2300 0.7600 2.8100 0.8800 ;
        RECT  2.5700 1.2950 2.8700 1.4150 ;
        RECT  0.2300 1.2700 2.6900 1.3900 ;
        RECT  1.8500 0.7100 2.0900 0.8800 ;
        RECT  1.9100 1.2700 2.0300 2.2100 ;
        RECT  1.0100 0.7100 1.2500 0.8800 ;
        RECT  1.0700 1.2700 1.1900 2.2100 ;
        RECT  0.3600 0.7600 0.5100 1.1450 ;
        RECT  0.3600 0.7600 0.4800 1.3900 ;
        RECT  0.2300 1.2700 0.3500 2.2100 ;
        RECT  0.2300 0.6400 0.3500 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  4.0100 -0.1800 4.1300 0.7050 ;
        RECT  3.1700 -0.1800 3.2900 0.7050 ;
        RECT  2.3300 -0.1800 2.4500 0.6400 ;
        RECT  1.4900 -0.1800 1.6100 0.6400 ;
        RECT  0.6500 -0.1800 0.7700 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  4.0100 1.4650 4.1300 2.7900 ;
        RECT  3.1700 1.4650 3.2900 2.7900 ;
        RECT  2.3300 1.5100 2.4500 2.7900 ;
        RECT  1.4900 1.5100 1.6100 2.7900 ;
        RECT  0.6500 1.5100 0.7700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.7100 2.1150 3.5900 2.1150 3.5900 1.1500 3.1900 1.1500 3.1900 1.1750 2.9500 1.1750
                 2.9500 1.1500 0.8700 1.1500 0.8700 1.0300 3.5900 1.0300 3.5900 0.6550 3.7100 0.6550 ;
    END
END BUFX8

MACRO BUFX6
    CLASS CORE ;
    FOREIGN BUFX6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8900 1.3900 2.0100 2.2100 ;
        RECT  0.1500 0.9100 2.0100 1.0300 ;
        RECT  1.8900 0.4000 2.0100 1.0300 ;
        RECT  0.2100 1.3900 2.0100 1.5100 ;
        RECT  1.0500 1.3900 1.1700 2.2100 ;
        RECT  0.9900 0.4000 1.1100 1.0300 ;
        RECT  0.3600 1.1750 0.5100 1.5100 ;
        RECT  0.3600 0.9100 0.4800 1.5100 ;
        RECT  0.2100 1.3900 0.3300 2.2100 ;
        RECT  0.1500 0.4000 0.2700 1.0300 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.8250 3.1200 1.2850 ;
        RECT  2.9700 0.8250 3.0900 1.3100 ;
        END
    END A
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  3.1500 1.4300 3.2700 2.7900 ;
        RECT  2.3100 1.4300 2.4300 2.7900 ;
        RECT  1.4700 1.6300 1.5900 2.7900 ;
        RECT  0.6300 1.6300 0.7500 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  3.1500 -0.1800 3.2700 0.7050 ;
        RECT  2.3100 -0.1800 2.4300 0.8950 ;
        RECT  1.4100 -0.1800 1.5300 0.7900 ;
        RECT  0.5700 -0.1800 0.6900 0.7900 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  2.8500 2.0800 2.7300 2.0800 2.7300 1.2700 0.7700 1.2700 0.7700 1.1500 2.7300 1.1500
                 2.7300 0.6550 2.8500 0.6550 ;
    END
END BUFX6

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9550 1.2400 2.0750 1.4800 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.8400 1.3600 2.0750 1.4800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3350 0.7100 1.5750 0.8300 ;
        RECT  1.3950 1.3200 1.5150 2.2100 ;
        RECT  0.5150 0.7600 1.4550 0.8800 ;
        RECT  0.5150 1.3200 1.5150 1.4400 ;
        RECT  0.5550 1.3200 0.8000 1.7250 ;
        RECT  0.5550 1.3200 0.6750 2.2100 ;
        RECT  0.5550 0.6400 0.6750 0.8800 ;
        RECT  0.5150 0.7600 0.6350 1.4400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.8150 -0.1800 1.9350 0.7000 ;
        RECT  0.9150 0.5200 1.1550 0.6400 ;
        RECT  0.9150 -0.1800 1.0350 0.6400 ;
        RECT  0.1350 -0.1800 0.2550 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8150 1.8450 1.9350 2.7900 ;
        RECT  0.9750 1.5600 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3550 2.2100 2.2350 2.2100 2.2350 1.1200 1.4150 1.1200 1.4150 1.1700 1.1750 1.1700
                 1.1750 1.1200 0.9950 1.1200 0.9950 1.1700 0.7550 1.1700 0.7550 1.0500 0.8750 1.0500
                 0.8750 1.0000 2.2350 1.0000 2.2350 0.6500 2.3550 0.6500 ;
    END
END BUFX4

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.0000 1.6700 1.5000 ;
        RECT  1.5200 1.0000 1.6700 1.4700 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6480  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9750 1.3200 1.0950 2.2100 ;
        RECT  0.9750 0.4000 1.0950 0.6400 ;
        RECT  0.1350 0.7600 1.0900 0.8800 ;
        RECT  0.1350 1.3200 1.0950 1.4400 ;
        RECT  0.9700 0.5200 1.0900 0.8800 ;
        RECT  0.3600 1.1750 0.5100 1.4400 ;
        RECT  0.3600 0.7600 0.4800 1.4400 ;
        RECT  0.1350 1.3200 0.2550 2.2100 ;
        RECT  0.1350 0.5900 0.2550 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3950 -0.1800 1.5150 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.3950 1.6200 1.5150 2.7900 ;
        RECT  0.5550 1.5600 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 2.2100 1.8150 2.2100 1.8150 0.8800 1.3300 0.8800 1.3300 1.1700 1.2100 1.1700
                 1.2100 0.7600 1.8150 0.7600 1.8150 0.5900 1.9350 0.5900 ;
    END
END BUFX3

MACRO BUFX20
    CLASS CORE ;
    FOREIGN BUFX20 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.8600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.5400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0200 1.2600 8.6200 1.3800 ;
        RECT  8.1350 1.2300 8.3950 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.6387  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9600 1.4250 7.0800 2.2100 ;
        RECT  0.3600 0.9450 7.0800 1.0650 ;
        RECT  6.9600 0.4000 7.0800 1.0650 ;
        RECT  0.2400 1.4250 7.0800 1.5450 ;
        RECT  6.1200 1.4250 6.2400 2.2100 ;
        RECT  6.1200 0.4000 6.2400 1.0650 ;
        RECT  5.2800 1.4250 5.4000 2.2100 ;
        RECT  5.2200 0.4000 5.3400 1.0650 ;
        RECT  4.4400 1.4250 4.5600 2.2100 ;
        RECT  4.3800 0.4000 4.5000 1.0650 ;
        RECT  3.6000 1.4250 3.7200 2.2100 ;
        RECT  3.5400 0.4000 3.6600 1.0650 ;
        RECT  2.7600 1.4250 2.8800 2.2100 ;
        RECT  2.7000 0.4000 2.8200 1.0650 ;
        RECT  1.9200 1.4250 2.0400 2.2100 ;
        RECT  1.8600 0.4000 1.9800 1.0650 ;
        RECT  1.0800 1.4250 1.2000 2.2100 ;
        RECT  1.0200 0.4000 1.1400 1.0650 ;
        RECT  0.3600 0.9450 0.5100 1.5450 ;
        RECT  0.3600 0.7850 0.4800 1.5450 ;
        RECT  0.2400 1.4250 0.3600 2.2100 ;
        RECT  0.1800 0.7850 0.4800 0.9050 ;
        RECT  0.1800 0.4000 0.3000 0.9050 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.8600 0.1800 ;
        RECT  9.0600 -0.1800 9.1800 0.7200 ;
        RECT  8.2200 -0.1800 8.3400 0.7200 ;
        RECT  7.3800 -0.1800 7.5000 0.9100 ;
        RECT  6.5400 -0.1800 6.6600 0.8250 ;
        RECT  5.6400 -0.1800 5.7600 0.8250 ;
        RECT  4.8000 -0.1800 4.9200 0.8250 ;
        RECT  3.9600 -0.1800 4.0800 0.8250 ;
        RECT  3.1200 -0.1800 3.2400 0.8250 ;
        RECT  2.2800 -0.1800 2.4000 0.8250 ;
        RECT  1.4400 -0.1800 1.5600 0.8250 ;
        RECT  0.6000 -0.1800 0.7200 0.8250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.8600 2.7900 ;
        RECT  9.0600 1.7400 9.1800 2.7900 ;
        RECT  8.2200 1.7400 8.3400 2.7900 ;
        RECT  7.3800 1.5600 7.5000 2.7900 ;
        RECT  6.5400 1.6650 6.6600 2.7900 ;
        RECT  5.7000 1.6650 5.8200 2.7900 ;
        RECT  4.8600 1.6650 4.9800 2.7900 ;
        RECT  4.0200 1.6650 4.1400 2.7900 ;
        RECT  3.1800 1.6650 3.3000 2.7900 ;
        RECT  2.3400 1.6650 2.4600 2.7900 ;
        RECT  1.5000 1.6650 1.6200 2.7900 ;
        RECT  0.6600 1.6650 0.7800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.6000 0.9600 7.9000 0.9600 7.9000 1.5000 9.6000 1.5000 9.6000 2.2100 9.4800 2.2100
                 9.4800 1.6200 8.7600 1.6200 8.7600 2.2100 8.6400 2.2100 8.6400 1.6200 7.9200 1.6200
                 7.9200 2.2100 7.8000 2.2100 7.8000 1.6200 7.7800 1.6200 7.7800 1.3050 0.8200 1.3050
                 0.8200 1.1850 7.7800 1.1850 7.7800 0.8400 7.8000 0.8400 7.8000 0.6700 7.9200 0.6700
                 7.9200 0.8400 8.6400 0.8400 8.6400 0.6700 8.7600 0.6700 8.7600 0.8400 9.4800 0.8400
                 9.4800 0.6700 9.6000 0.6700 ;
    END
END BUFX20

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2250 1.2750 1.3800 ;
        RECT  1.1550 1.1300 1.2750 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.2250 0.6750 2.1200 ;
        RECT  0.5550 0.6050 0.6750 0.8450 ;
        RECT  0.5150 0.7250 0.6350 1.3450 ;
        RECT  0.3600 0.8850 0.6350 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9750 -0.1800 1.0950 0.7700 ;
        RECT  0.1350 -0.1800 0.2550 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.5000 1.0950 2.7900 ;
        RECT  0.1350 1.4700 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5150 1.7400 1.3950 1.7400 1.3950 1.0100 1.0350 1.0100 1.0350 1.1050 0.7550 1.1050
                 0.7550 0.9850 0.9150 0.9850 0.9150 0.8900 1.3950 0.8900 1.3950 0.5300 1.5150 0.5300 ;
    END
END BUFX2

MACRO BUFX16
    CLASS CORE ;
    FOREIGN BUFX16 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.6850 1.2600 7.2850 1.3800 ;
        RECT  6.6850 1.2300 6.9450 1.3800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.7648  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5650 0.7150 5.8050 0.8350 ;
        RECT  5.6250 1.2950 5.7450 2.2100 ;
        RECT  0.5450 0.7650 5.6850 0.8850 ;
        RECT  0.5450 1.2950 5.7450 1.4150 ;
        RECT  4.7250 0.7150 4.9650 0.8850 ;
        RECT  4.7850 1.2950 4.9050 2.2100 ;
        RECT  3.8850 0.7150 4.1250 0.8850 ;
        RECT  3.9450 1.2950 4.0650 2.2100 ;
        RECT  3.0450 0.7150 3.2850 0.8850 ;
        RECT  3.1050 1.2950 3.2250 2.2100 ;
        RECT  2.2050 0.7150 2.4450 0.8850 ;
        RECT  2.2650 1.2950 2.3850 2.2100 ;
        RECT  1.3650 0.7150 1.6050 0.8850 ;
        RECT  1.4250 1.2950 1.5450 2.2100 ;
        RECT  0.5850 1.2950 0.8000 1.7250 ;
        RECT  0.5850 1.2950 0.7050 2.2100 ;
        RECT  0.5850 0.6450 0.7050 0.8850 ;
        RECT  0.5450 0.7650 0.6650 1.4150 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.7250 -0.1800 7.8450 0.7050 ;
        RECT  6.8850 -0.1800 7.0050 0.7050 ;
        RECT  6.0450 -0.1800 6.1650 0.7050 ;
        RECT  5.2050 -0.1800 5.3250 0.6450 ;
        RECT  4.3650 -0.1800 4.4850 0.6450 ;
        RECT  3.5250 -0.1800 3.6450 0.6450 ;
        RECT  2.6850 -0.1800 2.8050 0.6450 ;
        RECT  1.8450 -0.1800 1.9650 0.6450 ;
        RECT  1.0050 -0.1800 1.1250 0.6400 ;
        RECT  0.1650 -0.1800 0.2850 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.7250 1.5600 7.8450 2.7900 ;
        RECT  6.8850 1.7400 7.0050 2.7900 ;
        RECT  6.0450 1.5600 6.1650 2.7900 ;
        RECT  5.2050 1.5350 5.3250 2.7900 ;
        RECT  4.3650 1.5350 4.4850 2.7900 ;
        RECT  3.5250 1.5350 3.6450 2.7900 ;
        RECT  2.6850 1.5350 2.8050 2.7900 ;
        RECT  1.8450 1.5350 1.9650 2.7900 ;
        RECT  1.0050 1.5350 1.1250 2.7900 ;
        RECT  0.1650 1.4650 0.2850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.4250 0.9450 6.5650 0.9450 6.5650 1.5000 7.4250 1.5000 7.4250 2.2100 7.3050 2.2100
                 7.3050 1.6200 6.5850 1.6200 6.5850 2.2100 6.4650 2.2100 6.4650 1.6200 6.4450 1.6200
                 6.4450 1.1750 0.7850 1.1750 0.7850 1.0550 6.4450 1.0550 6.4450 0.8250 6.4650 0.8250
                 6.4650 0.6550 6.5850 0.6550 6.5850 0.8250 7.3050 0.8250 7.3050 0.6550 7.4250 0.6550 ;
    END
END BUFX16

MACRO BUFX12
    CLASS CORE ;
    FOREIGN BUFX12 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3240  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4500 1.3000 4.7750 1.4200 ;
        RECT  4.4200 1.4650 4.5700 1.7250 ;
        RECT  4.4500 1.3000 4.5700 1.7250 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.0736  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9150 1.3200 4.0350 2.2100 ;
        RECT  0.5150 0.8200 4.0350 0.9400 ;
        RECT  3.9150 0.4000 4.0350 0.9400 ;
        RECT  0.5150 1.3200 4.0350 1.4400 ;
        RECT  3.0750 1.3200 3.1950 2.2100 ;
        RECT  3.0750 0.4000 3.1950 0.9400 ;
        RECT  2.2350 1.3200 2.3550 2.2100 ;
        RECT  2.2350 0.4000 2.3550 0.9400 ;
        RECT  1.3950 1.3200 1.5150 2.2100 ;
        RECT  1.3950 0.4000 1.5150 0.9400 ;
        RECT  0.5550 1.3200 0.8000 1.7250 ;
        RECT  0.5550 1.3200 0.6750 2.2100 ;
        RECT  0.5550 0.4000 0.6750 0.9400 ;
        RECT  0.5150 0.8000 0.6350 1.4400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.1750 -0.1800 5.2950 0.7250 ;
        RECT  4.3350 -0.1800 4.4550 0.9150 ;
        RECT  3.4950 -0.1800 3.6150 0.7000 ;
        RECT  2.6550 -0.1800 2.7750 0.7000 ;
        RECT  1.8150 -0.1800 1.9350 0.7000 ;
        RECT  0.9750 -0.1800 1.0950 0.7000 ;
        RECT  0.1350 -0.1800 0.2550 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.1750 1.5600 5.2950 2.7900 ;
        RECT  4.3350 1.8450 4.4550 2.7900 ;
        RECT  3.4950 1.5600 3.6150 2.7900 ;
        RECT  2.6550 1.5600 2.7750 2.7900 ;
        RECT  1.8150 1.5600 1.9350 2.7900 ;
        RECT  0.9750 1.5600 1.0950 2.7900 ;
        RECT  0.1350 1.4300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7150 0.9650 5.0150 0.9650 5.0150 1.3200 5.7150 1.3200 5.7150 2.2100 5.5950 2.2100
                 5.5950 1.4400 5.0150 1.4400 5.0150 1.6600 4.8750 1.6600 4.8750 2.2100 4.7550 2.2100
                 4.7550 1.5400 4.8950 1.5400 4.8950 1.1800 3.9350 1.1800 3.9350 1.1950 3.6950 1.1950
                 3.6950 1.1800 3.0950 1.1800 3.0950 1.1950 2.8550 1.1950 2.8550 1.1800 2.6750 1.1800
                 2.6750 1.1950 2.4350 1.1950 2.4350 1.1800 1.8350 1.1800 1.8350 1.1950 1.5950 1.1950
                 1.5950 1.1800 0.9950 1.1800 0.9950 1.2000 0.7550 1.2000 0.7550 1.0800 0.8750 1.0800
                 0.8750 1.0600 4.7550 1.0600 4.7550 0.6750 4.8750 0.6750 4.8750 0.8450 5.5950 0.8450
                 5.5950 0.6750 5.7150 0.6750 ;
    END
END BUFX12

MACRO BMXIX4
    CLASS CORE ;
    FOREIGN BMXIX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN X2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0450 2.1100 6.3650 2.2500 ;
        RECT  6.1050 2.1000 6.3650 2.2500 ;
        RECT  5.5150 2.1100 6.3650 2.2300 ;
        RECT  5.5150 0.9500 5.6350 2.2300 ;
        RECT  5.0450 0.9500 5.6350 1.1900 ;
        END
    END X2
    PIN PPN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.3150 0.6800 8.4350 2.0100 ;
        RECT  7.4750 1.0250 8.4350 1.1450 ;
        RECT  7.4750 0.8850 7.7600 1.1450 ;
        RECT  7.4750 0.6800 7.5950 2.0100 ;
        END
    END PPN
    PIN M0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9900 2.0500 1.6200 2.1700 ;
        RECT  0.9900 1.6400 1.1100 2.1700 ;
        RECT  0.7250 1.6400 1.1100 1.7600 ;
        RECT  0.5600 1.5200 0.8550 1.6400 ;
        RECT  0.5950 1.6400 1.1100 1.6700 ;
        RECT  0.5600 1.1900 0.6800 1.6400 ;
        RECT  0.5200 1.1900 0.6800 1.4300 ;
        END
    END M0
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7400 2.0500 3.5600 2.1700 ;
        RECT  1.7400 1.8100 1.8600 2.1700 ;
        RECT  1.2300 1.8100 1.8600 1.9300 ;
        RECT  1.2300 1.4650 1.3800 1.9300 ;
        RECT  1.2300 1.2300 1.3500 1.9300 ;
        RECT  0.8000 1.2300 1.3500 1.3500 ;
        END
    END S
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 0.9950 2.2500 1.4500 ;
        RECT  2.1300 0.9800 2.2500 1.4500 ;
        END
    END A
    PIN M1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9600 1.3000 4.0800 1.4200 ;
        RECT  3.9600 1.1700 4.0800 1.4200 ;
        RECT  2.9150 1.2300 3.1750 1.3800 ;
        RECT  2.9600 0.3600 3.0800 1.4300 ;
        RECT  2.4600 0.3600 3.0800 0.4800 ;
        END
    END M1
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.7350 -0.1800 8.8550 0.7300 ;
        RECT  7.8950 -0.1800 8.0150 0.7300 ;
        RECT  7.0550 -0.1800 7.1750 0.9200 ;
        RECT  3.8800 -0.1800 4.0000 0.3800 ;
        RECT  2.0200 -0.1800 2.1400 0.8600 ;
        RECT  0.6800 -0.1800 0.8000 0.8300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  8.7350 1.3600 8.8550 2.7900 ;
        RECT  7.8950 1.3600 8.0150 2.7900 ;
        RECT  6.9950 2.0000 7.1150 2.7900 ;
        RECT  3.6600 2.2900 3.9000 2.7900 ;
        RECT  2.2400 2.2900 2.4800 2.7900 ;
        RECT  0.8400 2.2900 1.0800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.3150 1.8400 6.6700 1.8400 6.6700 1.9800 5.8750 1.9800 5.8750 1.9900 5.7550 1.9900
                 5.7550 0.8300 5.1450 0.8300 5.1450 0.6600 5.3850 0.6600 5.3850 0.7100 5.8750 0.7100
                 5.8750 1.8600 6.5500 1.8600 6.5500 1.7200 7.1950 1.7200 7.1950 1.0400 7.3150 1.0400 ;
        POLYGON  6.7550 1.6000 6.6350 1.6000 6.6350 0.9800 6.2350 0.9800 6.2350 0.8600 6.6350 0.8600
                 6.6350 0.6800 6.7550 0.6800 ;
        POLYGON  6.4250 1.7400 6.1850 1.7400 6.1850 1.5200 5.9950 1.5200 5.9950 0.5900 5.5650 0.5900
                 5.5650 0.4800 4.6650 0.4800 4.6650 1.9300 3.9200 1.9300 3.9200 1.6900 2.6750 1.6900
                 2.6750 0.8000 2.6000 0.8000 2.6000 0.6800 2.8400 0.6800 2.8400 0.8000 2.7950 0.8000
                 2.7950 1.5700 4.0400 1.5700 4.0400 1.8100 4.5450 1.8100 4.5450 0.3600 5.6850 0.3600
                 5.6850 0.4700 6.1150 0.4700 6.1150 1.4000 6.4250 1.4000 ;
        POLYGON  5.3950 2.1700 3.6800 2.1700 3.6800 1.9300 1.9800 1.9300 1.9800 1.6900 1.5000 1.6900
                 1.5000 0.7700 1.2600 0.7700 1.2600 0.6500 1.6200 0.6500 1.6200 1.5700 2.1000 1.5700
                 2.1000 1.8100 3.8000 1.8100 3.8000 2.0500 5.2750 2.0500 5.2750 1.4600 4.8050 1.4600
                 4.8050 0.8400 4.7850 0.8400 4.7850 0.6000 4.9050 0.6000 4.9050 0.7200 4.9250 0.7200
                 4.9250 1.3400 5.3950 1.3400 ;
        POLYGON  4.4250 0.9000 4.3200 0.9000 4.3200 1.5700 4.4000 1.5700 4.4000 1.6900 4.1600 1.6900
                 4.1600 1.5700 4.2000 1.5700 4.2000 1.0500 3.4400 1.0500 3.4400 1.1800 3.3200 1.1800
                 3.3200 0.9300 4.2000 0.9300 4.2000 0.7800 4.3050 0.7800 4.3050 0.6600 4.4250 0.6600 ;
        POLYGON  1.8600 1.4300 1.7400 1.4300 1.7400 0.5300 1.1400 0.5300 1.1400 0.9900 1.3600 0.9900
                 1.3600 1.1100 1.0200 1.1100 1.0200 1.0700 0.4000 1.0700 0.4000 1.5500 0.4400 1.5500
                 0.4400 1.7900 0.3200 1.7900 0.3200 1.6700 0.2800 1.6700 0.2800 0.9500 0.2600 0.9500
                 0.2600 0.5900 0.3800 0.5900 0.3800 0.8300 0.4000 0.8300 0.4000 0.9500 1.0200 0.9500
                 1.0200 0.4100 1.8600 0.4100 ;
    END
END BMXIX4

MACRO BMXIX2
    CLASS CORE ;
    FOREIGN BMXIX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN M0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2150 1.2300 1.3350 1.4900 ;
        RECT  0.3050 1.2300 1.3350 1.3500 ;
        RECT  0.3050 1.2300 0.5650 1.3800 ;
        RECT  0.3550 1.2300 0.4750 1.4700 ;
        END
    END M0
    PIN S
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7850 2.1100 3.4350 2.2300 ;
        RECT  1.0000 2.0300 2.9050 2.1500 ;
        RECT  1.0000 1.6100 1.1200 2.1500 ;
        RECT  0.7350 1.6100 1.1200 1.7300 ;
        RECT  0.5950 1.5200 0.9750 1.6700 ;
        RECT  0.7350 1.4700 0.9750 1.7300 ;
        END
    END S
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0450 1.1800 2.3050 1.3800 ;
        RECT  1.9550 1.2550 2.1950 1.4300 ;
        END
    END A
    PIN M1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7550 1.2500 3.9950 1.3700 ;
        RECT  2.9750 1.3100 3.8750 1.4300 ;
        RECT  3.2050 1.2300 3.4650 1.4300 ;
        END
    END M1
    PIN X2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1600 0.8850 6.3100 1.1450 ;
        RECT  6.1000 1.0250 6.2200 1.4500 ;
        END
    END X2
    PIN PPN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7850 0.6700 6.9050 1.0250 ;
        RECT  6.7800 0.8850 6.9000 1.9900 ;
        RECT  6.7400 0.8850 6.9000 1.1450 ;
        END
    END PPN
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  7.2050 -0.1800 7.3250 0.7200 ;
        RECT  6.2450 -0.1800 6.4850 0.3700 ;
        RECT  3.5550 -0.1800 3.7950 0.3200 ;
        RECT  1.9350 -0.1800 2.0550 0.8500 ;
        RECT  0.5550 -0.1800 0.6750 0.8500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  7.2000 1.3400 7.3200 2.7900 ;
        RECT  6.3600 1.5300 6.4800 2.7900 ;
        RECT  3.5550 2.2900 3.7950 2.7900 ;
        RECT  1.9950 2.2700 2.2350 2.7900 ;
        RECT  0.7150 1.8500 0.8350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.6200 1.2300 6.5000 1.2300 6.5000 0.6100 5.7050 0.6100 5.7050 0.5100 5.1350 0.5100
                 5.1350 1.7700 5.0150 1.7700 5.0150 0.3900 5.8250 0.3900 5.8250 0.4900 6.6200 0.4900 ;
        POLYGON  6.1200 1.7100 5.7950 1.7100 5.7950 2.2500 4.8750 2.2500 4.8750 2.1300 5.6750 2.1300
                 5.6750 1.2300 5.4950 1.2300 5.4950 0.9900 5.7650 0.9900 5.7650 0.7300 6.0050 0.7300
                 6.0050 0.8500 5.8850 0.8500 5.8850 1.1100 5.7950 1.1100 5.7950 1.5900 6.1200 1.5900 ;
        POLYGON  5.5550 0.8700 5.3750 0.8700 5.3750 1.6500 5.5550 1.6500 5.5550 2.0100 4.7550 2.0100
                 4.7550 2.1700 3.5550 2.1700 3.5550 1.9900 3.0250 1.9900 3.0250 1.9100 2.6950 1.9100
                 2.6950 1.7900 3.1450 1.7900 3.1450 1.8700 3.6750 1.8700 3.6750 2.0500 4.6350 2.0500
                 4.6350 1.8900 4.7750 1.8900 4.7750 0.5100 4.4150 0.5100 4.4150 0.5600 3.3000 0.5600
                 3.3000 0.6100 3.0350 0.6100 3.0350 0.8500 2.9150 0.8500 2.9150 0.4900 3.1800 0.4900
                 3.1800 0.4400 4.2950 0.4400 4.2950 0.3900 4.8950 0.3900 4.8950 1.8900 5.4350 1.8900
                 5.4350 1.7700 5.2550 1.7700 5.2550 0.7500 5.4350 0.7500 5.4350 0.6300 5.5550 0.6300 ;
        POLYGON  4.6550 0.8700 4.5150 0.8700 4.5150 1.5300 4.6550 1.5300 4.6550 1.7700 4.5150 1.7700
                 4.5150 1.9300 3.7950 1.9300 3.7950 1.6700 1.5750 1.6700 1.5750 1.9100 1.2950 1.9100
                 1.2950 1.7900 1.4550 1.7900 1.4550 0.7900 1.1350 0.7900 1.1350 0.6700 1.5750 0.6700
                 1.5750 1.5500 3.9150 1.5500 3.9150 1.8100 4.3950 1.8100 4.3950 0.7500 4.5350 0.7500
                 4.5350 0.6300 4.6550 0.6300 ;
        POLYGON  4.2750 0.8000 4.2350 0.8000 4.2350 1.5700 4.2750 1.5700 4.2750 1.6900 4.0350 1.6900
                 4.0350 1.5700 4.1150 1.5700 4.1150 1.1100 2.6150 1.1100 2.6150 1.4100 2.4950 1.4100
                 2.4950 0.9900 4.1150 0.9900 4.1150 0.8000 4.0350 0.8000 4.0350 0.6800 4.2750 0.6800 ;
        POLYGON  1.8150 1.4100 1.6950 1.4100 1.6950 0.5500 1.0150 0.5500 1.0150 0.9900 1.2350 0.9900
                 1.2350 1.1100 0.8950 1.1100 0.8950 1.0900 0.1850 1.0900 0.1850 1.7300 0.4150 1.7300
                 0.4150 1.9700 0.2950 1.9700 0.2950 1.8500 0.0650 1.8500 0.0650 0.7300 0.1350 0.7300
                 0.1350 0.6100 0.2550 0.6100 0.2550 0.9700 0.8950 0.9700 0.8950 0.4300 1.8150 0.4300 ;
    END
END BMXIX2

MACRO AOI33XL
    CLASS CORE ;
    FOREIGN AOI33XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 0.8500 1.6700 1.2250 ;
        RECT  1.5450 0.8500 1.6650 1.4850 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8050 1.0400 0.9250 1.2950 ;
        RECT  0.6500 1.0400 0.9250 1.1600 ;
        RECT  0.6500 0.8850 0.8000 1.1600 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.8800 2.5400 1.3500 ;
        RECT  2.3900 0.8500 2.5100 1.3500 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8750 0.8500 2.0850 1.1000 ;
        RECT  1.7900 0.8750 2.0250 1.1450 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.8500 1.3800 1.2200 ;
        RECT  1.2250 1.1000 1.3450 1.4750 ;
        END
    END A2
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.7950 0.5100 1.4300 ;
        RECT  0.3600 0.7950 0.5100 1.1700 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2928  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6600 1.4650 2.8300 1.7250 ;
        RECT  2.6600 0.6100 2.7800 1.7250 ;
        RECT  2.6450 1.4700 2.7650 1.8300 ;
        RECT  1.3850 0.6100 2.7800 0.7300 ;
        RECT  1.8050 1.4700 2.8300 1.5900 ;
        RECT  1.8050 1.4700 1.9250 1.8300 ;
        RECT  1.3850 0.4000 1.5050 0.7300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  2.4450 0.3700 2.6850 0.4900 ;
        RECT  2.4450 -0.1800 2.5650 0.4900 ;
        RECT  0.3250 -0.1800 0.4450 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  0.9050 2.2300 1.0250 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3450 1.9500 2.1650 1.9500 2.1650 2.0700 1.3850 2.0700 1.3850 1.8300 0.4850 1.8300
                 0.4850 1.7100 1.5050 1.7100 1.5050 1.9500 2.0450 1.9500 2.0450 1.8300 2.2250 1.8300
                 2.2250 1.7100 2.3450 1.7100 ;
    END
END AOI33XL

MACRO AOI33X4
    CLASS CORE ;
    FOREIGN AOI33X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.7300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.8550 0.7500 9.9750 1.1700 ;
        RECT  5.3750 0.7500 9.9750 0.8700 ;
        RECT  7.5000 0.7500 7.7400 1.0900 ;
        RECT  5.2350 0.9400 5.4950 1.0900 ;
        RECT  5.3750 0.7500 5.4950 1.0900 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7550 0.7500 4.8750 1.1500 ;
        RECT  4.7100 0.7500 4.8750 1.1450 ;
        RECT  0.5750 0.7500 4.8750 0.8700 ;
        RECT  2.6400 0.7500 2.8800 1.0900 ;
        RECT  0.5750 0.7500 0.6950 1.1500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2900 0.9900 4.5900 1.1100 ;
        RECT  2.4000 1.2100 3.4350 1.3300 ;
        RECT  3.2900 0.9900 3.4350 1.3300 ;
        RECT  2.4000 1.0600 2.5200 1.3300 ;
        RECT  1.3400 1.0600 2.5200 1.1800 ;
        RECT  0.8550 1.1750 1.4600 1.2950 ;
        RECT  1.2300 1.1750 1.3800 1.4350 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.3500 1.1750 9.6550 1.3800 ;
        RECT  9.5350 1.1400 9.6550 1.3800 ;
        RECT  9.3500 1.1750 9.5000 1.4350 ;
        RECT  9.0100 1.1750 9.6550 1.2950 ;
        RECT  9.0100 1.0400 9.1300 1.2950 ;
        RECT  7.8600 1.0400 9.1300 1.1600 ;
        RECT  7.0650 1.2100 7.9800 1.3300 ;
        RECT  7.8600 1.0400 7.9800 1.3300 ;
        RECT  7.0650 0.9900 7.1850 1.3300 ;
        RECT  5.7950 0.9900 7.1850 1.1100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.6350 1.2800 8.8750 1.4000 ;
        RECT  6.7800 1.4500 8.7550 1.5700 ;
        RECT  8.6350 1.2800 8.7550 1.5700 ;
        RECT  6.7800 1.2300 6.9450 1.5700 ;
        RECT  6.6350 1.2800 6.9450 1.4000 ;
        RECT  6.6850 1.2300 6.9450 1.4000 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.2300 4.0450 1.3800 ;
        RECT  2.1600 1.4500 3.8700 1.5700 ;
        RECT  3.7500 1.2600 3.9050 1.4800 ;
        RECT  2.1600 1.3000 2.2800 1.5700 ;
        RECT  1.6150 1.3000 2.2800 1.4200 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.7984  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.7950 1.5600 9.9150 2.0100 ;
        RECT  5.5950 1.6900 9.9150 1.8100 ;
        RECT  8.9550 1.5600 9.0750 2.0100 ;
        RECT  1.5350 0.5100 8.9350 0.6300 ;
        RECT  8.1150 1.6900 8.2350 2.0100 ;
        RECT  7.2750 1.6900 7.3950 2.0100 ;
        RECT  6.4350 1.5600 6.5550 2.0100 ;
        RECT  5.5950 1.2300 5.7150 2.0100 ;
        RECT  4.9950 1.2300 5.7150 1.3800 ;
        RECT  4.9950 1.1800 5.1500 1.4300 ;
        RECT  4.9950 0.5100 5.1150 1.4300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.7300 0.1800 ;
        RECT  9.9550 0.4600 10.1950 0.5800 ;
        RECT  9.9550 -0.1800 10.0750 0.5800 ;
        RECT  7.6750 -0.1800 7.9150 0.3900 ;
        RECT  5.0350 -0.1800 5.2750 0.3900 ;
        RECT  2.5550 -0.1800 2.7950 0.3900 ;
        RECT  0.3750 0.4600 0.6150 0.5800 ;
        RECT  0.3750 -0.1800 0.4950 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.7300 2.7900 ;
        RECT  4.7550 1.9300 4.8750 2.7900 ;
        RECT  3.9150 1.9300 4.0350 2.7900 ;
        RECT  3.0750 1.9300 3.1950 2.7900 ;
        RECT  2.2350 1.9300 2.3550 2.7900 ;
        RECT  1.3950 1.9300 1.5150 2.7900 ;
        RECT  0.5550 1.9300 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.3350 2.2500 5.1750 2.2500 5.1750 1.8100 4.4550 1.8100 4.4550 2.2100 4.3350 2.2100
                 4.3350 1.8100 3.6150 1.8100 3.6150 2.2100 3.4950 2.2100 3.4950 1.8100 2.7750 1.8100
                 2.7750 2.2100 2.6550 2.2100 2.6550 1.8100 1.9350 1.8100 1.9350 2.2100 1.8150 2.2100
                 1.8150 1.8100 1.0950 1.8100 1.0950 2.2100 0.9750 2.2100 0.9750 1.8100 0.2550 1.8100
                 0.2550 2.2100 0.1350 2.2100 0.1350 1.5600 0.2550 1.5600 0.2550 1.6900 0.9750 1.6900
                 0.9750 1.5600 1.0950 1.5600 1.0950 1.6900 1.8150 1.6900 1.8150 1.5600 1.9350 1.5600
                 1.9350 1.6900 4.3350 1.6900 4.3350 1.5600 4.4550 1.5600 4.4550 1.6900 5.1750 1.6900
                 5.1750 1.5600 5.2950 1.5600 5.2950 2.1300 6.0150 2.1300 6.0150 1.9300 6.1350 1.9300
                 6.1350 2.1300 6.8550 2.1300 6.8550 1.9300 6.9750 1.9300 6.9750 2.1300 7.6950 2.1300
                 7.6950 1.9300 7.8150 1.9300 7.8150 2.1300 8.5350 2.1300 8.5350 1.9300 8.6550 1.9300
                 8.6550 2.1300 9.3750 2.1300 9.3750 1.9300 9.4950 1.9300 9.4950 2.1300 10.2150 2.1300
                 10.2150 1.5600 10.3350 1.5600 ;
    END
END AOI33X4

MACRO AOI33X2
    CLASS CORE ;
    FOREIGN AOI33X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8150 0.7500 4.9350 1.1700 ;
        RECT  3.0000 0.7500 4.9350 0.8700 ;
        RECT  3.0000 0.7500 3.1200 1.1700 ;
        RECT  2.9700 0.8850 3.1200 1.1450 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.3900 0.7500 2.5100 1.1700 ;
        RECT  0.4750 0.7500 2.5100 0.8700 ;
        RECT  0.4750 0.7500 0.5950 1.1500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7550 0.9900 2.2500 1.1100 ;
        RECT  0.9400 0.9900 1.0900 1.4350 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4200 0.9900 4.6150 1.2300 ;
        RECT  4.4200 0.9900 4.5700 1.4350 ;
        RECT  3.2750 0.9900 4.6150 1.1100 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4950 1.2300 3.8350 1.4400 ;
        RECT  3.4950 1.2300 3.7550 1.4650 ;
        END
    END B2
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.2300 1.8850 1.4350 ;
        RECT  1.4650 1.2300 1.7700 1.4600 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.8992  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7550 1.5600 4.8750 2.0100 ;
        RECT  3.0750 1.5850 4.8750 1.7050 ;
        RECT  3.9150 1.5600 4.0350 2.0100 ;
        RECT  1.5300 0.5100 3.9950 0.6300 ;
        RECT  3.0750 1.5500 3.1950 2.0100 ;
        RECT  2.6250 1.5500 3.1950 1.6700 ;
        RECT  2.6250 1.5200 2.8850 1.6700 ;
        RECT  2.7300 0.5100 2.8500 1.6700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.9150 0.4600 5.1550 0.5800 ;
        RECT  4.9150 -0.1800 5.0350 0.5800 ;
        RECT  2.6500 -0.1800 2.8900 0.3900 ;
        RECT  0.2750 0.4600 0.5150 0.5800 ;
        RECT  0.2750 -0.1800 0.3950 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  2.1750 2.0300 2.4150 2.1500 ;
        RECT  2.1750 2.0300 2.2950 2.7900 ;
        RECT  1.3350 2.0300 1.5750 2.1500 ;
        RECT  1.3350 2.0300 1.4550 2.7900 ;
        RECT  0.4950 2.0300 0.7350 2.1500 ;
        RECT  0.4950 2.0300 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.2950 2.2500 2.6550 2.2500 2.6550 1.9100 1.9350 1.9100 1.9350 2.2100 1.8150 2.2100
                 1.8150 1.9100 1.0950 1.9100 1.0950 2.2100 0.9750 2.2100 0.9750 1.9100 0.2550 1.9100
                 0.2550 2.2100 0.1350 2.2100 0.1350 1.5600 0.2550 1.5600 0.2550 1.7900 0.9750 1.7900
                 0.9750 1.5600 1.0950 1.5600 1.0950 1.7900 1.8150 1.7900 1.8150 1.5800 1.9350 1.5800
                 1.9350 1.7900 2.7750 1.7900 2.7750 2.1300 3.4950 2.1300 3.4950 1.8250 3.6150 1.8250
                 3.6150 2.1300 4.3350 2.1300 4.3350 1.8250 4.4550 1.8250 4.4550 2.1300 5.1750 2.1300
                 5.1750 1.5600 5.2950 1.5600 ;
    END
END AOI33X2

MACRO AOI33X1
    CLASS CORE ;
    FOREIGN AOI33X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5700 1.0300 1.6900 1.4550 ;
        RECT  1.5200 1.0300 1.6900 1.4350 ;
        END
    END B2
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 0.8850 1.0900 1.1850 ;
        RECT  0.8500 0.8800 0.9700 1.1700 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0000 2.5400 1.4700 ;
        RECT  2.3900 1.0000 2.5100 1.5000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1750 2.1300 1.2950 ;
        RECT  2.0100 1.0550 2.1300 1.2950 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.0000 1.3800 1.4550 ;
        RECT  1.2300 1.0000 1.3500 1.4850 ;
        END
    END A2
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.7600 0.5100 1.2350 ;
        RECT  0.3600 0.7600 0.5100 1.2150 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.5276  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.4650 2.8300 1.7250 ;
        RECT  2.6900 1.4650 2.8100 2.2100 ;
        RECT  2.6800 0.7600 2.8000 1.7400 ;
        RECT  1.8500 1.6200 2.8100 1.7400 ;
        RECT  1.4300 0.7600 2.8000 0.8800 ;
        RECT  1.8500 1.5600 1.9700 2.0100 ;
        RECT  1.4300 0.5900 1.5500 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.4900 -0.1800 2.6100 0.6400 ;
        RECT  0.3700 -0.1800 0.4900 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  1.0100 1.8450 1.1300 2.7900 ;
        RECT  0.1700 1.5600 0.2900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3900 2.2500 1.4300 2.2500 1.4300 1.7250 0.7100 1.7250 0.7100 2.2100 0.5900 2.2100
                 0.5900 1.5600 0.7100 1.5600 0.7100 1.6050 1.5500 1.6050 1.5500 2.1300 2.2700 2.1300
                 2.2700 1.8600 2.3900 1.8600 ;
    END
END AOI33X1

MACRO AOI32XL
    CLASS CORE ;
    FOREIGN AOI32XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7750 0.5100 1.2350 ;
        RECT  0.3800 0.7750 0.5000 1.2650 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1750 0.9950 2.2950 1.4350 ;
        RECT  2.1000 0.7750 2.2500 1.1950 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0400 0.7250 1.1600 1.0550 ;
        RECT  0.9400 0.5950 1.0900 0.9300 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6550 0.6150 1.7750 1.0550 ;
        RECT  1.5200 0.7750 1.6700 1.1950 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.7350 0.8200 1.1050 ;
        RECT  0.6500 0.4900 0.8000 0.8550 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2388  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9350 1.3150 2.0550 1.6750 ;
        RECT  1.2300 1.3150 2.0550 1.4350 ;
        RECT  1.3200 0.4150 1.4400 0.6550 ;
        RECT  1.2300 1.1750 1.4000 1.4350 ;
        RECT  1.2800 0.5350 1.4000 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  2.1550 -0.1800 2.2750 0.6550 ;
        RECT  0.2200 -0.1800 0.3400 0.6550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.0950 2.0750 1.2150 2.7900 ;
        RECT  0.1350 2.0750 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4750 1.7950 2.2950 1.7950 2.2950 1.9150 1.5150 1.9150 1.5150 1.6750 0.5550 1.6750
                 0.5550 1.5550 1.6350 1.5550 1.6350 1.7950 2.1750 1.7950 2.1750 1.6750 2.3550 1.6750
                 2.3550 1.5550 2.4750 1.5550 ;
    END
END AOI32XL

MACRO AOI32X4
    CLASS CORE ;
    FOREIGN AOI32X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.9900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.5250 0.9900 8.5250 1.1100 ;
        RECT  5.5250 0.9400 5.7850 1.1100 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9250 0.9900 5.1650 1.1100 ;
        RECT  5.0000 0.8850 5.1500 1.1450 ;
        RECT  5.0000 0.7500 5.1200 1.1450 ;
        RECT  0.7450 0.7500 5.1200 0.8700 ;
        RECT  2.9050 0.7500 3.1450 1.0900 ;
        RECT  0.7450 0.7500 0.8650 1.1500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4600 1.0000 4.8050 1.1200 ;
        RECT  2.6650 1.2100 3.5800 1.3300 ;
        RECT  3.4600 1.0000 3.5800 1.3300 ;
        RECT  2.6650 1.0600 2.7850 1.3300 ;
        RECT  2.1350 1.0600 2.7850 1.1800 ;
        RECT  1.0250 0.9900 2.2550 1.1100 ;
        RECT  1.2300 0.9900 1.3800 1.4350 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.1850 1.2600 7.7850 1.3800 ;
        RECT  6.3950 1.2300 6.6550 1.3800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4250 1.4500 3.9250 1.5700 ;
        RECT  3.8050 1.2400 3.9250 1.5700 ;
        RECT  2.4250 1.3000 2.5450 1.5700 ;
        RECT  1.7850 1.3000 2.5450 1.4200 ;
        RECT  1.7550 1.2300 2.0150 1.3800 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2850 1.5000 8.4050 2.0100 ;
        RECT  5.7650 1.5000 8.4050 1.6200 ;
        RECT  1.7050 0.5100 7.6650 0.6300 ;
        RECT  7.4450 1.5000 7.5650 2.0100 ;
        RECT  6.6050 1.5000 6.7250 2.0100 ;
        RECT  5.7650 1.3200 5.8850 2.0100 ;
        RECT  5.2850 1.2300 5.7850 1.4400 ;
        RECT  5.2850 0.5100 5.4050 1.4400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.9900 0.1800 ;
        RECT  8.1250 -0.1800 8.2450 0.6400 ;
        RECT  6.7250 -0.1800 6.9650 0.3900 ;
        RECT  5.2450 -0.1800 5.4850 0.3900 ;
        RECT  2.7250 -0.1800 2.9650 0.3900 ;
        RECT  0.5450 0.4600 0.7850 0.5800 ;
        RECT  0.5450 -0.1800 0.6650 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.9900 2.7900 ;
        RECT  4.9250 1.9300 5.0450 2.7900 ;
        RECT  4.0850 1.9300 4.2050 2.7900 ;
        RECT  3.2450 1.9300 3.3650 2.7900 ;
        RECT  2.4050 1.9300 2.5250 2.7900 ;
        RECT  1.5650 1.9300 1.6850 2.7900 ;
        RECT  0.7250 1.9300 0.8450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.8250 2.2500 5.3450 2.2500 5.3450 1.8100 4.6250 1.8100 4.6250 2.2100 4.5050 2.2100
                 4.5050 1.8100 3.7850 1.8100 3.7850 2.2100 3.6650 2.2100 3.6650 1.8100 2.9450 1.8100
                 2.9450 2.2100 2.8250 2.2100 2.8250 1.8100 2.1050 1.8100 2.1050 2.2100 1.9850 2.2100
                 1.9850 1.8100 1.2650 1.8100 1.2650 2.2100 1.1450 2.2100 1.1450 1.8100 0.4250 1.8100
                 0.4250 2.2100 0.3050 2.2100 0.3050 1.5600 0.4250 1.5600 0.4250 1.6900 1.1450 1.6900
                 1.1450 1.5600 1.2650 1.5600 1.2650 1.6900 1.9850 1.6900 1.9850 1.5600 2.1050 1.5600
                 2.1050 1.6900 4.5050 1.6900 4.5050 1.5600 4.6250 1.5600 4.6250 1.6900 5.3450 1.6900
                 5.3450 1.5600 5.4650 1.5600 5.4650 2.1300 6.1850 2.1300 6.1850 1.7400 6.3050 1.7400
                 6.3050 2.1300 7.0250 2.1300 7.0250 1.7400 7.1450 1.7400 7.1450 2.1300 7.8650 2.1300
                 7.8650 1.7400 7.9850 1.7400 7.9850 2.1300 8.7050 2.1300 8.7050 1.5600 8.8250 1.5600 ;
    END
END AOI32X4

MACRO AOI32X2
    CLASS CORE ;
    FOREIGN AOI32X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1100 0.9900 4.3500 1.1100 ;
        RECT  3.2050 0.9350 4.2300 1.0550 ;
        RECT  3.0050 0.9900 3.4650 1.0900 ;
        RECT  3.0050 0.9900 3.3250 1.1100 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4200 0.8200 2.5400 1.1500 ;
        RECT  2.3900 0.8200 2.5400 1.1450 ;
        RECT  0.5250 0.8200 2.5400 0.9400 ;
        RECT  0.5250 0.8200 0.6450 1.1500 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7050 1.1950 3.9900 1.4350 ;
        RECT  3.8400 1.1750 3.9900 1.4350 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  0.8050 1.0600 2.2200 1.1800 ;
        RECT  2.0800 1.1750 2.2500 1.3000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3150 1.3000 1.5550 1.4200 ;
        RECT  1.1750 1.5200 1.4350 1.6700 ;
        RECT  1.3150 1.3000 1.4350 1.6700 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9650 1.5550 4.0850 2.0100 ;
        RECT  3.1250 1.5550 4.0850 1.6750 ;
        RECT  1.5400 0.5800 3.7250 0.7000 ;
        RECT  3.1250 1.5200 3.2450 2.0100 ;
        RECT  2.6250 1.5200 3.2450 1.6400 ;
        RECT  2.6250 1.5200 2.8850 1.6700 ;
        RECT  2.7650 0.5800 2.8850 1.6700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  4.1850 -0.1800 4.3050 0.6400 ;
        RECT  2.6850 0.3400 2.9250 0.4600 ;
        RECT  2.6850 -0.1800 2.8050 0.4600 ;
        RECT  0.3250 0.4600 0.5650 0.5800 ;
        RECT  0.3250 -0.1800 0.4450 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  2.2250 2.0300 2.4650 2.1500 ;
        RECT  2.2250 2.0300 2.3450 2.7900 ;
        RECT  1.3850 2.0300 1.6250 2.1500 ;
        RECT  1.3850 2.0300 1.5050 2.7900 ;
        RECT  0.5450 2.0300 0.7850 2.1500 ;
        RECT  0.5450 2.0300 0.6650 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.5050 2.2500 2.7050 2.2500 2.7050 1.9100 1.9850 1.9100 1.9850 2.2100 1.8650 2.2100
                 1.8650 1.9100 1.1450 1.9100 1.1450 2.2100 1.0250 2.2100 1.0250 1.9100 0.3050 1.9100
                 0.3050 2.2100 0.1850 2.2100 0.1850 1.5600 0.3050 1.5600 0.3050 1.7900 1.8650 1.7900
                 1.8650 1.5600 1.9850 1.5600 1.9850 1.7900 2.8250 1.7900 2.8250 2.1300 3.5450 2.1300
                 3.5450 1.7950 3.6650 1.7950 3.6650 2.1300 4.3850 2.1300 4.3850 1.5600 4.5050 1.5600 ;
    END
END AOI32X2

MACRO AOI32X1
    CLASS CORE ;
    FOREIGN AOI32X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7800 0.5100 1.2150 ;
        RECT  0.3800 0.7800 0.5000 1.3200 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1350 1.0250 2.5400 1.1450 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.1350 1.0250 2.2550 1.2650 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0400 0.8200 1.1600 1.1700 ;
        RECT  0.9400 0.5950 1.0900 0.9450 ;
        END
    END A2
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9400 2.0150 1.0950 ;
        RECT  1.5200 0.9850 1.8750 1.1100 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.8450 0.8200 1.2700 ;
        RECT  0.6500 0.5600 0.8000 0.9650 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3778  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8150 1.2600 1.9350 2.0100 ;
        RECT  1.2800 1.2600 1.9350 1.3800 ;
        RECT  1.2800 1.2300 1.7250 1.3800 ;
        RECT  1.3200 0.6100 1.4400 0.8650 ;
        RECT  1.2800 0.7450 1.4000 1.3800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  2.0800 -0.1800 2.2000 0.6600 ;
        RECT  0.2200 -0.1800 0.3400 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.5000 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3550 2.2500 1.3950 2.2500 1.3950 1.6200 0.6750 1.6200 0.6750 2.1500 0.5550 2.1500
                 0.5550 1.5000 1.5150 1.5000 1.5150 2.1300 2.2350 2.1300 2.2350 1.5000 2.3550 1.5000 ;
    END
END AOI32X1

MACRO AOI31XL
    CLASS CORE ;
    FOREIGN AOI31XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.6600 0.8200 1.1050 ;
        RECT  0.6500 0.7200 0.8000 1.1450 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1150 0.8850 1.2350 1.2450 ;
        RECT  0.9400 0.8850 1.2350 1.2400 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8150 1.1250 1.9350 1.5200 ;
        RECT  1.4650 1.1550 1.9350 1.3800 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.2900 0.8850 0.5300 1.0900 ;
        RECT  0.3600 0.8850 0.5100 1.2800 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1992  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.0550 1.1750 2.2500 1.4350 ;
        RECT  2.0550 0.8850 2.1750 1.6850 ;
        RECT  1.3750 0.8850 2.1750 1.0050 ;
        RECT  1.3750 0.5250 1.4950 1.0050 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.7950 -0.1800 1.9150 0.7650 ;
        RECT  0.2200 -0.1800 0.3400 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.0950 2.0850 1.2150 2.7900 ;
        RECT  0.1350 2.0850 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6950 1.7450 1.5750 1.7450 1.5750 1.6250 0.5550 1.6250 0.5550 1.5050 1.6950 1.5050 ;
    END
END AOI31XL

MACRO AOI31X4
    CLASS CORE ;
    FOREIGN AOI31X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6550 1.2300 5.2500 1.3500 ;
        RECT  4.6550 1.2300 4.9150 1.3800 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.3300 1.2250 6.9100 1.3450 ;
        RECT  6.3950 1.2250 6.6550 1.3800 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3100 1.2600 3.5500 1.3800 ;
        RECT  2.6250 1.2300 3.4300 1.3500 ;
        RECT  2.6250 1.2300 2.8850 1.3800 ;
        RECT  2.6250 1.0100 2.8500 1.3800 ;
        RECT  2.6100 1.0100 2.8500 1.1300 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0500 1.2600 1.8700 1.3800 ;
        RECT  1.0500 1.2300 1.4350 1.3800 ;
        RECT  1.0500 1.0100 1.1700 1.3800 ;
        RECT  0.9300 1.0100 1.1700 1.1300 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0696  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.4000 0.6800 7.5200 0.9200 ;
        RECT  7.2200 0.8000 7.5200 0.9200 ;
        RECT  4.0400 0.8500 7.3400 0.9700 ;
        RECT  7.0300 1.4650 7.1800 1.7250 ;
        RECT  7.0300 0.8500 7.1500 1.7250 ;
        RECT  7.0100 1.5000 7.1300 2.0100 ;
        RECT  6.1700 1.5000 7.1800 1.6200 ;
        RECT  6.5600 0.6800 6.6800 0.9700 ;
        RECT  6.1700 1.5000 6.2900 2.0100 ;
        RECT  5.7200 0.6800 5.8400 0.9700 ;
        RECT  4.8800 0.6800 5.0000 0.9700 ;
        RECT  4.0400 0.6800 4.1600 0.9700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  6.9800 -0.1800 7.1000 0.7300 ;
        RECT  6.1400 -0.1800 6.2600 0.7300 ;
        RECT  1.5500 -0.1800 1.6700 0.6500 ;
        RECT  0.7100 -0.1800 0.8300 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  5.3300 1.7400 5.4500 2.7900 ;
        RECT  4.4900 1.7400 4.6100 2.7900 ;
        RECT  3.6500 1.7400 3.7700 2.7900 ;
        RECT  2.8100 1.7400 2.9300 2.7900 ;
        RECT  1.9700 1.7400 2.0900 2.7900 ;
        RECT  1.1300 1.7400 1.2500 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.5500 2.2500 5.7500 2.2500 5.7500 1.6200 5.0300 1.6200 5.0300 2.2100 4.9100 2.2100
                 4.9100 1.6200 4.1900 1.6200 4.1900 2.2100 4.0700 2.2100 4.0700 1.6200 3.3500 1.6200
                 3.3500 2.2100 3.2300 2.2100 3.2300 1.6200 2.5100 1.6200 2.5100 2.2100 2.3900 2.2100
                 2.3900 1.6200 1.6700 1.6200 1.6700 2.2100 1.5500 2.2100 1.5500 1.6200 0.8300 1.6200
                 0.8300 2.2100 0.7100 2.2100 0.7100 1.5000 5.8700 1.5000 5.8700 2.1300 6.5900 2.1300
                 6.5900 1.7400 6.7100 1.7400 6.7100 2.1300 7.4300 2.1300 7.4300 1.5600 7.5500 1.5600 ;
        POLYGON  5.4200 0.7300 5.3000 0.7300 5.3000 0.4800 4.5800 0.4800 4.5800 0.7300 4.4600 0.7300
                 4.4600 0.4800 3.3500 0.4800 3.3500 0.6500 3.2300 0.6500 3.2300 0.4800 2.5100 0.4800
                 2.5100 0.6500 2.3900 0.6500 2.3900 0.3600 5.4200 0.3600 ;
        POLYGON  3.7700 0.8900 0.2900 0.8900 0.2900 0.6000 0.4100 0.6000 0.4100 0.7700 1.1300 0.7700
                 1.1300 0.6000 1.2500 0.6000 1.2500 0.7700 1.9700 0.7700 1.9700 0.6000 2.0900 0.6000
                 2.0900 0.7700 2.8100 0.7700 2.8100 0.6000 2.9300 0.6000 2.9300 0.7700 3.6500 0.7700
                 3.6500 0.6000 3.7700 0.6000 ;
    END
END AOI31X4

MACRO AOI31X2
    CLASS CORE ;
    FOREIGN AOI31X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 0.7600 3.4100 1.2100 ;
        RECT  3.2600 0.7600 3.3800 1.2350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3200 0.8850 2.5400 1.1450 ;
        RECT  2.3200 0.7500 2.5100 1.1450 ;
        RECT  2.3200 0.7500 2.4400 1.1500 ;
        RECT  0.4800 0.7500 2.5100 0.8700 ;
        RECT  0.4800 0.7500 0.6000 1.1500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7600 0.9900 2.1600 1.1100 ;
        RECT  0.9400 0.9900 1.0900 1.4350 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.2300 1.7250 1.5000 ;
        END
    END A2
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0800 1.3550 3.2000 2.0100 ;
        RECT  2.9700 1.1750 3.1200 1.4350 ;
        RECT  3.0000 0.4000 3.1200 1.4750 ;
        RECT  1.4400 0.5100 3.1200 0.6300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.4200 -0.1800 3.5400 0.6400 ;
        RECT  2.4600 -0.1800 2.7000 0.3900 ;
        RECT  0.2800 0.4600 0.5200 0.5800 ;
        RECT  0.2800 -0.1800 0.4000 0.5800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  2.2400 1.8600 2.3600 2.7900 ;
        RECT  1.4000 1.8600 1.5200 2.7900 ;
        RECT  0.5600 1.8600 0.6800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.6200 2.2500 2.6600 2.2500 2.6600 1.7400 1.9400 1.7400 1.9400 2.2100 1.8200 2.2100
                 1.8200 1.7400 1.1000 1.7400 1.1000 2.2100 0.9800 2.2100 0.9800 1.7400 0.2600 1.7400
                 0.2600 2.2100 0.1400 2.2100 0.1400 1.5600 0.2600 1.5600 0.2600 1.6200 0.9800 1.6200
                 0.9800 1.5600 1.1000 1.5600 1.1000 1.6200 2.6600 1.6200 2.6600 1.5600 2.7800 1.5600
                 2.7800 2.1300 3.5000 2.1300 3.5000 1.5600 3.6200 1.5600 ;
    END
END AOI31X2

MACRO AOI31X1
    CLASS CORE ;
    FOREIGN AOI31X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8150 1.0050 0.9350 1.2500 ;
        RECT  0.6500 1.0050 0.9350 1.1450 ;
        RECT  0.6500 0.8800 0.8000 1.1450 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 1.0000 1.3800 1.4350 ;
        RECT  1.2100 1.0000 1.3300 1.4600 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5500 1.0000 1.6700 1.4750 ;
        RECT  1.5200 1.0000 1.6700 1.4500 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.9700 0.5100 1.4400 ;
        RECT  0.3900 0.9400 0.5100 1.4400 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3196  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.8850 1.9600 1.1450 ;
        RECT  1.8150 0.7600 1.9350 2.2100 ;
        RECT  1.8100 0.7600 1.9350 1.1450 ;
        RECT  1.2950 0.7600 1.9350 0.8800 ;
        RECT  1.2950 0.5900 1.4150 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.7150 -0.1800 1.8350 0.6400 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  0.9750 1.8200 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5150 2.2100 1.3950 2.2100 1.3950 1.7150 1.2150 1.7150 1.2150 1.7000 0.6750 1.7000
                 0.6750 2.2100 0.5550 2.2100 0.5550 1.5600 0.6750 1.5600 0.6750 1.5800 1.3350 1.5800
                 1.3350 1.5950 1.5150 1.5950 ;
    END
END AOI31X1

MACRO AOI2BB2XL
    CLASS CORE ;
    FOREIGN AOI2BB2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1920  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5450 1.5300 2.7850 1.6500 ;
        RECT  2.5650 0.7000 2.6850 1.6500 ;
        RECT  1.5500 0.7000 2.6850 0.8200 ;
        RECT  1.5200 0.8850 1.6700 1.1450 ;
        RECT  1.5500 0.7000 1.6700 1.1450 ;
        END
    END Y
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.2650 0.5100 1.7300 ;
        RECT  0.3600 1.2350 0.4800 1.7300 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 0.8500 0.8550 1.2200 ;
        RECT  0.5950 0.9050 0.8550 1.1150 ;
        END
    END A0N
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2550 0.9700 2.4450 1.2100 ;
        RECT  2.0000 0.9400 2.3750 1.0900 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.8850 1.1500 3.1750 1.3800 ;
        RECT  2.8850 1.0000 3.0050 1.4100 ;
        END
    END B0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.8250 -0.1800 2.9450 0.8800 ;
        RECT  1.4250 -0.1800 1.6650 0.3400 ;
        RECT  0.5550 -0.1800 0.6750 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  1.7650 1.5800 1.8850 2.7900 ;
        RECT  0.5950 1.9700 0.7150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.2050 1.7600 3.0850 1.7600 3.0850 1.8900 2.3050 1.8900 2.3050 1.6400 2.0050 1.6400
                 2.0050 1.4600 1.4650 1.4600 1.4650 1.7000 1.3450 1.7000 1.3450 1.3400 2.1250 1.3400
                 2.1250 1.5200 2.4250 1.5200 2.4250 1.7700 2.9650 1.7700 2.9650 1.6400 3.2050 1.6400 ;
        POLYGON  2.2050 0.4800 2.0850 0.4800 2.0850 0.5800 0.9150 0.5800 0.9150 0.6600 0.2550 0.6600
                 0.2550 0.9000 0.2400 0.9000 0.2400 1.8500 0.2950 1.8500 0.2950 2.0900 0.1750 2.0900
                 0.1750 1.9700 0.1200 1.9700 0.1200 0.7800 0.1350 0.7800 0.1350 0.5400 0.7950 0.5400
                 0.7950 0.4600 1.9650 0.4600 1.9650 0.3600 2.2050 0.3600 ;
        POLYGON  1.4000 1.2200 1.2800 1.2200 1.2800 1.1000 1.1550 1.1000 1.1550 2.0900 1.1350 2.0900
                 1.1350 2.2100 1.0150 2.2100 1.0150 1.9700 1.0350 1.9700 1.0350 0.7200 1.2750 0.7200
                 1.2750 0.8400 1.1550 0.8400 1.1550 0.9800 1.4000 0.9800 ;
    END
END AOI2BB2XL

MACRO AOI2BB2X4
    CLASS CORE ;
    FOREIGN AOI2BB2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0100 0.5100 1.4800 ;
        RECT  0.3750 1.0100 0.4950 1.5100 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0100 0.8350 1.3900 ;
        RECT  0.6500 1.0650 0.8000 1.4350 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3650 0.9900 7.8250 1.1100 ;
        RECT  7.3650 0.4100 7.4850 1.1100 ;
        RECT  6.5650 0.4100 7.4850 0.5300 ;
        RECT  6.5650 0.4100 6.6850 1.0900 ;
        RECT  4.9450 0.9700 6.6850 1.0900 ;
        RECT  4.9450 0.9400 5.2050 1.0900 ;
        RECT  4.9250 0.9900 5.1650 1.1100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6850 1.2600 7.0050 1.3800 ;
        RECT  5.8150 1.2300 6.0750 1.3800 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5850 1.5000 7.7050 2.0100 ;
        RECT  4.9450 1.5000 7.7050 1.6200 ;
        RECT  7.1250 0.6500 7.2450 1.6200 ;
        RECT  6.9050 0.6500 7.2450 0.7700 ;
        RECT  6.7450 1.5000 6.8650 2.0100 ;
        RECT  5.9050 1.5000 6.0250 2.0100 ;
        RECT  5.1600 0.6500 5.6650 0.7700 ;
        RECT  2.8500 0.7000 5.2800 0.8200 ;
        RECT  4.9450 1.5000 5.2050 1.6700 ;
        RECT  5.0650 1.5000 5.1850 2.0100 ;
        RECT  4.9450 1.2300 5.0650 1.6700 ;
        RECT  4.6850 1.2300 5.0650 1.3500 ;
        RECT  4.6850 0.7000 4.8050 1.3500 ;
        RECT  3.7450 0.6500 3.9850 0.8200 ;
        RECT  2.4650 0.6500 2.9700 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  7.6050 -0.1800 7.7250 0.6400 ;
        RECT  6.3250 -0.1800 6.4450 0.6400 ;
        RECT  4.5850 0.4600 4.8250 0.5800 ;
        RECT  4.5850 -0.1800 4.7050 0.5800 ;
        RECT  3.1050 0.4600 3.3450 0.5800 ;
        RECT  3.1050 -0.1800 3.2250 0.5800 ;
        RECT  1.8850 -0.1800 2.0050 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.6500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  4.1650 1.7100 4.4050 2.1500 ;
        RECT  4.1650 1.7100 4.2850 2.7900 ;
        RECT  3.3850 1.7100 3.5050 2.7900 ;
        RECT  2.5450 1.7100 2.6650 2.7900 ;
        RECT  1.7050 1.7100 1.8250 2.7900 ;
        RECT  0.5550 1.6300 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  8.1250 2.2500 4.6450 2.2500 4.6450 1.5900 3.9250 1.5900 3.9250 2.2100 3.8050 2.2100
                 3.8050 1.5900 3.0850 1.5900 3.0850 2.2100 2.9650 2.2100 2.9650 1.5900 2.2450 1.5900
                 2.2450 2.2100 2.1250 2.2100 2.1250 1.5900 1.4050 1.5900 1.4050 2.2100 1.2850 2.2100
                 1.2850 1.4700 4.7650 1.4700 4.7650 2.1300 5.4850 2.1300 5.4850 1.7400 5.6050 1.7400
                 5.6050 2.1300 6.3250 2.1300 6.3250 1.7400 6.4450 1.7400 6.4450 2.1300 7.1650 2.1300
                 7.1650 1.7400 7.2850 1.7400 7.2850 2.1300 8.0050 2.1300 8.0050 1.5600 8.1250 1.5600 ;
        POLYGON  4.5650 1.3500 1.1550 1.3500 1.1550 1.6800 1.0950 1.6800 1.0950 1.8000 0.9750 1.8000
                 0.9750 1.5600 1.0350 1.5600 1.0350 0.6000 1.1550 0.6000 1.1550 1.2300 4.5650 1.2300 ;
        POLYGON  3.8250 1.1100 2.2250 1.1100 2.2250 0.8800 1.4300 0.8800 1.4300 0.4800 0.9150 0.4800
                 0.9150 0.8900 0.2400 0.8900 0.2400 1.6000 0.2550 1.6000 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.7200 0.1200 1.7200 0.1200 0.7200 0.1350 0.7200 0.1350 0.6000 0.2550 0.6000
                 0.2550 0.7700 0.7950 0.7700 0.7950 0.3600 1.5500 0.3600 1.5500 0.7600 2.3450 0.7600
                 2.3450 0.9900 3.8250 0.9900 ;
    END
END AOI2BB2X4

MACRO AOI2BB2X2
    CLASS CORE ;
    FOREIGN AOI2BB2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.9300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0800 0.5100 1.4350 ;
        RECT  0.3850 0.9000 0.5050 1.4350 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7250 0.9050 0.8450 1.2400 ;
        RECT  0.6500 0.8100 0.8000 1.1450 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2000 0.9900 4.4400 1.1100 ;
        RECT  3.4950 0.9700 4.3200 1.0900 ;
        RECT  3.4950 0.9400 3.7550 1.0900 ;
        RECT  3.2400 0.9900 3.6650 1.1100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7850 1.2100 4.0450 1.4250 ;
        RECT  3.6650 1.2300 4.0450 1.4200 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.2550 1.5450 4.3750 2.0100 ;
        RECT  3.0000 1.5450 4.3750 1.6650 ;
        RECT  3.2300 0.6500 3.9600 0.7700 ;
        RECT  3.4150 1.5450 3.5350 2.0100 ;
        RECT  2.2150 0.7300 3.3500 0.8500 ;
        RECT  3.0000 0.7300 3.1200 1.6650 ;
        RECT  2.9700 1.1750 3.1200 1.4350 ;
        RECT  2.0950 0.6500 2.3350 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.9300 0.1800 ;
        RECT  4.4200 -0.1800 4.5400 0.6400 ;
        RECT  2.8700 0.4600 3.1100 0.5800 ;
        RECT  2.8700 -0.1800 2.9900 0.5800 ;
        RECT  1.5150 -0.1800 1.6350 0.6400 ;
        RECT  0.5550 -0.1800 0.6750 0.4000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.9300 2.7900 ;
        RECT  2.5150 2.0250 2.7550 2.1500 ;
        RECT  2.5150 2.0250 2.6350 2.7900 ;
        RECT  1.7350 1.7100 1.8550 2.7900 ;
        RECT  0.6150 2.0150 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.7950 2.2100 4.7500 2.2100 4.7500 2.2500 3.0400 2.2500 3.0400 2.2100 2.9950 2.2100
                 2.9950 1.9050 2.4200 1.9050 2.4200 1.5900 2.2750 1.5900 2.2750 2.2100 2.1550 2.2100
                 2.1550 1.5900 1.4350 1.5900 1.4350 2.2100 1.3150 2.2100 1.3150 1.4700 2.5400 1.4700
                 2.5400 1.7850 3.1150 1.7850 3.1150 2.0900 3.1600 2.0900 3.1600 2.1300 3.8350 2.1300
                 3.8350 1.7850 3.9550 1.7850 3.9550 2.1300 4.6300 2.1300 4.6300 2.0900 4.6750 2.0900
                 4.6750 1.5600 4.7950 1.5600 ;
        POLYGON  2.8500 1.3500 1.1550 1.3500 1.1550 1.4700 1.1250 1.4700 1.1250 1.6150 1.0050 1.6150
                 1.0050 1.3500 1.0350 1.3500 1.0350 0.6800 1.1550 0.6800 1.1550 1.2300 2.8500 1.2300 ;
        POLYGON  2.1750 1.1100 1.8550 1.1100 1.8550 0.8800 1.2750 0.8800 1.2750 0.5600 0.9150 0.5600
                 0.9150 0.6800 0.2550 0.6800 0.2550 0.9200 0.2400 0.9200 0.2400 1.5550 0.3150 1.5550
                 0.3150 1.6750 0.0750 1.6750 0.0750 1.5550 0.1200 1.5550 0.1200 0.8000 0.1350 0.8000
                 0.1350 0.5600 0.7950 0.5600 0.7950 0.4400 1.3950 0.4400 1.3950 0.7600 1.9750 0.7600
                 1.9750 0.9900 2.1750 0.9900 ;
    END
END AOI2BB2X2

MACRO AOI2BB2X1
    CLASS CORE ;
    FOREIGN AOI2BB2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 0.7600 2.8000 2.0100 ;
        RECT  2.3900 0.7600 2.8000 0.8800 ;
        RECT  2.2000 0.6500 2.5400 0.7700 ;
        RECT  2.3900 0.5950 2.5400 0.8800 ;
        END
    END Y
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4400 1.0250 0.8000 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        RECT  0.4400 1.0250 0.5600 1.2650 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7600 1.2650 0.8800 1.5650 ;
        RECT  0.6500 1.4150 0.8000 1.7250 ;
        END
    END A0N
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0250 2.5400 1.4800 ;
        RECT  2.4200 1.0000 2.5400 1.4800 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.8850 3.1200 1.3550 ;
        RECT  2.9600 0.9000 3.0800 1.4000 ;
        END
    END B0
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.9000 -0.1800 3.0200 0.6400 ;
        RECT  1.6200 -0.1800 1.7400 0.6400 ;
        RECT  0.6600 -0.1800 0.7800 0.5250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  1.8400 1.8400 1.9600 2.7900 ;
        RECT  0.6000 1.8450 0.7200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.2200 2.2100 3.1750 2.2100 3.1750 2.2500 2.2600 2.2500 2.2600 1.7200 1.5400 1.7200
                 1.5400 2.2100 1.4200 2.2100 1.4200 1.5600 1.5400 1.5600 1.5400 1.6000 2.3800 1.6000
                 2.3800 2.1300 3.0550 2.1300 3.0550 2.0900 3.1000 2.0900 3.1000 1.5600 3.2200 1.5600 ;
        POLYGON  2.2200 1.1700 1.9600 1.1700 1.9600 0.8800 1.3800 0.8800 1.3800 0.4800 1.0200 0.4800
                 1.0200 0.7650 0.3000 0.7650 0.3000 1.9650 0.1800 1.9650 0.1800 0.6000 0.3000 0.6000
                 0.3000 0.6450 0.9000 0.6450 0.9000 0.3600 1.5000 0.3600 1.5000 0.7600 2.0800 0.7600
                 2.0800 0.9300 2.2200 0.9300 ;
        POLYGON  1.7600 1.3200 1.2600 1.3200 1.2600 1.8450 1.1400 1.8450 1.1400 1.9650 1.0200 1.9650
                 1.0200 1.7250 1.1400 1.7250 1.1400 0.6000 1.2600 0.6000 1.2600 1.2000 1.7600 1.2000 ;
    END
END AOI2BB2X1

MACRO AOI2BB1XL
    CLASS CORE ;
    FOREIGN AOI2BB1XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7500 0.8200 1.9600 1.1600 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 1.3150 1.3800 1.7250 ;
        RECT  1.2100 1.3000 1.3300 1.7250 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.4650 1.0100 1.6250 ;
        RECT  0.8900 1.3850 1.0100 1.6250 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1776  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5700 0.5200 0.8100 0.6400 ;
        RECT  0.2500 0.8200 0.6900 0.9400 ;
        RECT  0.5700 0.5200 0.6900 0.9400 ;
        RECT  0.4100 1.3000 0.5300 1.9650 ;
        RECT  0.0700 1.3000 0.5300 1.4200 ;
        RECT  0.0700 1.1750 0.3700 1.4200 ;
        RECT  0.2500 0.8200 0.3700 1.4200 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.8900 -0.1800 2.0100 0.7000 ;
        RECT  1.0500 -0.1800 1.1700 0.7000 ;
        RECT  0.2100 -0.1800 0.3300 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.0500 1.8450 1.1700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.8700 1.9050 1.5000 1.9050 1.5000 1.1800 0.4900 1.1800 0.4900 1.0600 1.5000 1.0600
                 1.5000 0.7000 1.4700 0.7000 1.4700 0.4600 1.5900 0.4600 1.5900 0.5800 1.6200 0.5800
                 1.6200 1.7850 1.8700 1.7850 ;
    END
END AOI2BB1XL

MACRO AOI2BB1X4
    CLASS CORE ;
    FOREIGN AOI2BB1X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4200 1.0400 3.3200 1.1600 ;
        RECT  0.6500 1.0400 0.8000 1.4350 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1300 0.9850 4.2800 1.4400 ;
        RECT  4.1300 0.9650 4.2500 1.4400 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5500 0.7800 3.7000 1.2350 ;
        RECT  3.5800 0.7600 3.7000 1.2350 ;
        END
    END A0N
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9664  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1800 0.7600 3.2000 0.8800 ;
        RECT  3.0800 0.5900 3.2000 0.8800 ;
        RECT  2.2600 1.5950 2.3800 2.2100 ;
        RECT  2.2400 0.5900 2.3600 0.8800 ;
        RECT  0.1800 1.5950 2.3800 1.7150 ;
        RECT  1.4000 0.5900 1.5200 0.8800 ;
        RECT  0.9800 1.5600 1.1000 2.2100 ;
        RECT  0.5600 0.5900 0.6800 0.8800 ;
        RECT  0.3050 1.5950 0.5650 1.9600 ;
        RECT  0.1800 1.5950 0.5650 1.9300 ;
        RECT  0.1800 0.7600 0.3000 1.9300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  4.3400 -0.1800 4.4600 0.6400 ;
        RECT  3.5000 -0.1800 3.6200 0.6400 ;
        RECT  2.6600 -0.1800 2.7800 0.6400 ;
        RECT  1.8200 -0.1800 1.9400 0.6400 ;
        RECT  0.9800 -0.1800 1.1000 0.6400 ;
        RECT  0.1400 -0.1800 0.2600 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  3.3000 1.5950 3.4200 2.7900 ;
        RECT  1.6200 1.8350 1.7400 2.7900 ;
        RECT  0.2200 2.0800 0.4600 2.2000 ;
        RECT  0.2200 2.0800 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.0600 2.2100 3.9400 2.2100 3.9400 1.6800 3.8900 1.6800 3.8900 1.4750 1.2200 1.4750
                 1.2200 1.4000 1.0800 1.4000 1.0800 1.2800 1.3400 1.2800 1.3400 1.3550 2.3200 1.3550
                 2.3200 1.3000 2.5600 1.3000 2.5600 1.3550 3.8900 1.3550 3.8900 0.7250 3.9200 0.7250
                 3.9200 0.5900 4.0400 0.5900 4.0400 0.8450 4.0100 0.8450 4.0100 1.5600 4.0600 1.5600 ;
    END
END AOI2BB1X4

MACRO AOI2BB1X2
    CLASS CORE ;
    FOREIGN AOI2BB1X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.0450 2.5400 1.5000 ;
        RECT  2.3900 1.0250 2.5100 1.5000 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8950 0.8300 2.0150 1.1950 ;
        RECT  1.8100 0.8050 1.9600 1.1650 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4150 1.0600 1.6350 1.1800 ;
        RECT  0.6500 1.0600 0.8000 1.4350 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1750 0.8050 1.5150 0.9250 ;
        RECT  1.3950 0.6350 1.5150 0.9250 ;
        RECT  0.9750 1.5550 1.0950 2.2100 ;
        RECT  0.1750 1.5550 1.0950 1.6750 ;
        RECT  0.5550 0.6350 0.6750 0.9250 ;
        RECT  0.1750 0.8050 0.2950 1.6750 ;
        RECT  0.0700 1.1750 0.2950 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.7150 -0.1800 2.8350 0.8750 ;
        RECT  1.8150 -0.1800 1.9350 0.6850 ;
        RECT  0.9750 -0.1800 1.0950 0.6850 ;
        RECT  0.1350 -0.1800 0.2550 0.6850 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  1.6150 1.5600 1.7350 2.7900 ;
        RECT  0.3350 1.7950 0.4550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.4950 1.7400 2.1500 1.7400 2.1500 1.4350 1.1750 1.4350 1.1750 1.4200 1.0550 1.4200
                 1.0550 1.3000 1.2950 1.3000 1.2950 1.3150 2.1500 1.3150 2.1500 0.7850 2.2950 0.7850
                 2.2950 0.6350 2.4150 0.6350 2.4150 0.9050 2.2700 0.9050 2.2700 1.6200 2.4950 1.6200 ;
    END
END AOI2BB1X2

MACRO AOI2BB1X1
    CLASS CORE ;
    FOREIGN AOI2BB1X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.0950 1.9600 1.4350 ;
        RECT  1.7800 0.9800 1.9000 1.3200 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.4100 1.3800 1.7250 ;
        RECT  1.2400 1.2200 1.3600 1.7250 ;
        END
    END A0N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6800 1.3400 0.9800 1.4600 ;
        RECT  0.8600 1.2200 0.9800 1.4600 ;
        RECT  0.6500 1.4650 0.8000 1.7250 ;
        RECT  0.6800 1.3400 0.8000 1.7250 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3196  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6000 0.6900 0.8400 0.8100 ;
        RECT  0.2400 0.7400 0.7200 0.8600 ;
        RECT  0.3800 1.2700 0.5000 2.2100 ;
        RECT  0.2400 1.2700 0.5000 1.3900 ;
        RECT  0.2400 0.7400 0.3600 1.3900 ;
        RECT  0.0700 0.8850 0.3600 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.9200 -0.1800 2.0400 0.8600 ;
        RECT  1.0800 -0.1800 1.2000 0.8600 ;
        RECT  0.1800 0.5000 0.4200 0.6200 ;
        RECT  0.1800 -0.1800 0.3000 0.6200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.0200 1.8450 1.1400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9000 1.7400 1.5000 1.7400 1.5000 1.1000 0.7400 1.1000 0.7400 1.1500 0.4800 1.1500
                 0.4800 1.0300 0.6200 1.0300 0.6200 0.9800 1.5000 0.9800 1.5000 0.6200 1.6200 0.6200
                 1.6200 1.6200 1.9000 1.6200 ;
    END
END AOI2BB1X1

MACRO AOI22XL
    CLASS CORE ;
    FOREIGN AOI22XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.6800 0.8200 1.0400 ;
        RECT  0.6500 0.5000 0.8000 0.8550 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 0.5000 1.3800 0.9600 ;
        RECT  1.2100 0.4700 1.3300 0.9600 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5700 0.8000 1.6900 1.2350 ;
        RECT  1.5200 0.8850 1.6700 1.3000 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7850 0.5100 1.2400 ;
        RECT  0.3600 0.7600 0.4800 1.2400 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1932  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.4800 1.5150 1.7200 ;
        RECT  1.2150 1.4800 1.5150 1.6000 ;
        RECT  1.2150 1.0800 1.3350 1.6000 ;
        RECT  0.9700 1.0800 1.3350 1.2000 ;
        RECT  0.9400 0.8850 1.0900 1.1450 ;
        RECT  0.9700 0.4000 1.0900 1.2000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.7100 -0.1800 1.8300 0.6400 ;
        RECT  0.2000 -0.1800 0.3200 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  0.5550 1.6000 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 1.8400 1.7550 1.8400 1.7550 1.9600 0.9750 1.9600 0.9750 1.4800 0.3150 1.4800
                 0.3150 1.6600 0.0750 1.6600 0.0750 1.5400 0.1950 1.5400 0.1950 1.3600 1.0950 1.3600
                 1.0950 1.8400 1.6350 1.8400 1.6350 1.7200 1.8150 1.7200 1.8150 1.6000 1.9350 1.6000 ;
    END
END AOI22XL

MACRO AOI22X4
    CLASS CORE ;
    FOREIGN AOI22X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.2500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7150 0.9900 6.6750 1.1100 ;
        RECT  3.7850 0.9400 4.0450 1.1100 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.9900 3.3550 1.1800 ;
        RECT  3.2350 0.9400 3.3550 1.1800 ;
        RECT  2.9700 0.9900 3.1200 1.4350 ;
        RECT  0.4350 0.9900 3.3550 1.1100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2550 1.2300 2.7750 1.3500 ;
        RECT  1.4650 1.2300 1.7250 1.3800 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3550 1.2600 5.8750 1.3800 ;
        RECT  5.5250 1.2300 5.7850 1.3800 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.3824  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4350 1.5000 6.5550 2.0100 ;
        RECT  3.9150 1.5000 6.5550 1.6200 ;
        RECT  5.5950 1.5000 5.7150 2.0100 ;
        RECT  5.4750 0.6500 5.7150 0.7700 ;
        RECT  1.5350 0.7000 5.5950 0.8200 ;
        RECT  4.7550 1.5000 4.8750 2.0100 ;
        RECT  4.1950 0.6500 4.4350 0.8200 ;
        RECT  3.9150 1.3150 4.0350 2.0100 ;
        RECT  3.4750 1.3150 4.0350 1.4350 ;
        RECT  3.4750 1.2300 3.7550 1.4350 ;
        RECT  3.4750 0.7000 3.5950 1.4350 ;
        RECT  2.6950 0.6500 2.9350 0.8200 ;
        RECT  1.4150 0.6500 1.6550 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.2500 0.1800 ;
        RECT  6.1750 -0.1800 6.2950 0.6400 ;
        RECT  4.8350 0.4600 5.0750 0.5800 ;
        RECT  4.8350 -0.1800 4.9550 0.5800 ;
        RECT  3.4350 0.4600 3.6750 0.5800 ;
        RECT  3.4350 -0.1800 3.5550 0.5800 ;
        RECT  2.0550 0.4600 2.2950 0.5800 ;
        RECT  2.0550 -0.1800 2.1750 0.5800 ;
        RECT  0.8350 -0.1800 0.9550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.2500 2.7900 ;
        RECT  3.0750 1.7950 3.1950 2.7900 ;
        RECT  2.2350 1.7950 2.3550 2.7900 ;
        RECT  1.3950 1.7950 1.5150 2.7900 ;
        RECT  0.5550 1.7950 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.9750 2.2500 3.4950 2.2500 3.4950 1.6750 2.7750 1.6750 2.7750 2.2100 2.6550 2.2100
                 2.6550 1.6750 1.9350 1.6750 1.9350 2.2100 1.8150 2.2100 1.8150 1.6750 1.0950 1.6750
                 1.0950 2.2100 0.9750 2.2100 0.9750 1.6750 0.2550 1.6750 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.5550 3.6150 1.5550 3.6150 2.1300 4.3350 2.1300 4.3350 1.7400 4.4550 1.7400
                 4.4550 2.1300 5.1750 2.1300 5.1750 1.7400 5.2950 1.7400 5.2950 2.1300 6.0150 2.1300
                 6.0150 1.7400 6.1350 1.7400 6.1350 2.1300 6.8550 2.1300 6.8550 1.5600 6.9750 1.5600 ;
    END
END AOI22X4

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5000 0.9900 1.7750 1.1100 ;
        RECT  0.5950 0.9400 1.6200 0.9900 ;
        RECT  0.7350 0.8700 1.6200 0.9900 ;
        RECT  0.5550 0.9700 0.8550 1.0900 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0950 0.9400 3.4650 1.0900 ;
        RECT  3.0950 0.9400 3.3350 1.1100 ;
        RECT  2.4400 0.8700 3.3250 0.9900 ;
        RECT  2.1350 0.9900 2.5600 1.1100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6800 1.1400 2.8300 1.6100 ;
        RECT  2.6800 1.1100 2.8000 1.6100 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.1100 1.3800 1.5800 ;
        RECT  1.2550 1.1100 1.3750 1.6100 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0950 1.5600 3.2150 2.0100 ;
        RECT  2.2550 1.7300 3.2150 1.8500 ;
        RECT  1.0550 0.6300 2.8550 0.7500 ;
        RECT  2.2550 1.2600 2.3750 2.0100 ;
        RECT  1.7550 1.2600 2.3750 1.3800 ;
        RECT  1.7550 1.2300 2.0150 1.3800 ;
        RECT  1.8950 0.6300 2.0150 1.3800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.3150 -0.1800 3.4350 0.6400 ;
        RECT  1.8350 0.3900 2.0750 0.5100 ;
        RECT  1.8350 -0.1800 1.9550 0.5100 ;
        RECT  0.4750 -0.1800 0.5950 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  1.4150 1.9700 1.5350 2.7900 ;
        RECT  0.5750 1.9700 0.6950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.6350 2.2500 1.8350 2.2500 1.8350 1.8500 1.1150 1.8500 1.1150 2.2100 0.9950 2.2100
                 0.9950 1.8500 0.2750 1.8500 0.2750 2.2100 0.1550 2.2100 0.1550 1.5600 0.2750 1.5600
                 0.2750 1.7300 0.9950 1.7300 0.9950 1.7000 1.1150 1.7000 1.1150 1.7300 1.8350 1.7300
                 1.8350 1.5600 1.9550 1.5600 1.9550 2.1300 2.6750 2.1300 2.6750 1.9700 2.7950 1.9700
                 2.7950 2.1300 3.5150 2.1300 3.5150 1.5600 3.6350 1.5600 ;
    END
END AOI22X2

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.7350 0.8200 1.1700 ;
        RECT  0.6500 0.5950 0.8000 1.0050 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 0.7950 1.3800 1.2150 ;
        RECT  1.2100 0.7950 1.3300 1.2350 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 0.7850 1.6700 1.2350 ;
        RECT  1.5300 0.7600 1.6500 1.2350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.8850 0.5100 1.3400 ;
        RECT  0.3800 0.8850 0.5000 1.3600 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3478  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.3550 1.5150 2.0100 ;
        RECT  0.9700 1.3550 1.5150 1.4750 ;
        RECT  0.9400 1.1750 1.0900 1.4350 ;
        RECT  0.9700 0.5900 1.0900 1.4750 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.6900 -0.1800 1.8100 0.6400 ;
        RECT  0.2200 -0.1800 0.3400 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  0.5550 1.8350 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9350 2.2500 0.9750 2.2500 0.9750 1.7150 0.2550 1.7150 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.5600 0.2550 1.5600 0.2550 1.5950 1.0950 1.5950 1.0950 2.1300 1.8150 2.1300
                 1.8150 1.5600 1.9350 1.5600 ;
    END
END AOI22X1

MACRO AOI222XL
    CLASS CORE ;
    FOREIGN AOI222XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 0.9150 1.1450 1.1050 ;
        RECT  0.7050 0.8800 1.0050 1.0350 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3700 0.7100 2.5400 1.1450 ;
        RECT  2.3700 0.7100 2.4900 1.1700 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4650 ;
        RECT  1.8750 1.3100 2.2500 1.4450 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3450 0.7600 0.5850 1.0000 ;
        RECT  0.3050 0.8300 0.5650 1.0900 ;
        END
    END A0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6100 1.2650 2.8500 1.3850 ;
        RECT  2.6800 0.8850 2.8300 1.1450 ;
        RECT  2.6800 0.8850 2.8000 1.3850 ;
        END
    END C1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 0.8250 1.7250 1.0900 ;
        RECT  1.4500 0.7600 1.6900 1.0050 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3384  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 0.8850 3.1200 1.1450 ;
        RECT  2.5150 1.5050 3.0900 1.6250 ;
        RECT  2.9700 0.4700 3.0900 1.6250 ;
        RECT  2.8500 0.4000 2.9700 0.6400 ;
        RECT  1.2550 0.4700 3.0900 0.5900 ;
        RECT  2.5150 1.5050 2.6350 1.8650 ;
        RECT  1.2550 0.4000 1.3750 0.6400 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  1.9900 -0.1800 2.2300 0.3500 ;
        RECT  0.2850 -0.1800 0.4050 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  0.9850 2.1350 1.1050 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.0550 1.9850 2.8750 1.9850 2.8750 2.1050 1.3150 2.1050 1.3150 1.9250 1.1950 1.9250
                 1.1950 1.8050 1.4350 1.8050 1.4350 1.9850 2.0950 1.9850 2.0950 1.7450 2.2150 1.7450
                 2.2150 1.9850 2.7550 1.9850 2.7550 1.8650 2.9350 1.8650 2.9350 1.7450 3.0550 1.7450 ;
        POLYGON  1.7950 1.8650 1.6750 1.8650 1.6750 1.6850 0.6250 1.6850 0.6250 1.8300 0.5050 1.8300
                 0.5050 1.5650 1.7950 1.5650 ;
    END
END AOI222XL

MACRO AOI222X4
    CLASS CORE ;
    FOREIGN AOI222X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 11.0200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2750 1.0200 3.5150 1.1400 ;
        RECT  0.5150 0.9900 3.3950 1.1100 ;
        RECT  1.9950 0.9900 2.2350 1.1400 ;
        RECT  0.5950 0.9400 0.8550 1.1100 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6250 0.9900 10.5050 1.1100 ;
        RECT  10.1650 0.9400 10.4250 1.1100 ;
        RECT  8.7850 0.9900 9.0250 1.1400 ;
        RECT  7.5050 1.0200 7.7450 1.1400 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.0050 1.0200 7.2450 1.1400 ;
        RECT  4.3650 0.9900 7.1250 1.1100 ;
        RECT  5.4550 0.9900 5.6950 1.1400 ;
        RECT  4.3650 1.2300 4.6250 1.3800 ;
        RECT  4.3650 0.9900 4.4850 1.3800 ;
        RECT  4.1650 1.0200 4.4850 1.1400 ;
        END
    END B0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.1450 1.2600 9.6650 1.3800 ;
        RECT  9.2950 1.2300 9.5550 1.3800 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3550 1.2600 2.8750 1.3800 ;
        RECT  1.4650 1.2300 1.7250 1.3800 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9050 1.2600 6.4050 1.3800 ;
        RECT  5.8150 1.2300 6.0750 1.3800 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.6576  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  10.2650 1.5000 10.3850 2.0100 ;
        RECT  3.9250 1.5000 10.3850 1.6200 ;
        RECT  9.4250 1.5000 9.5450 2.0100 ;
        RECT  9.2650 0.6800 9.5050 0.8000 ;
        RECT  1.6350 0.7300 9.3850 0.8500 ;
        RECT  8.5850 1.5000 8.7050 2.0100 ;
        RECT  7.9850 0.6800 8.2250 0.8500 ;
        RECT  7.7450 1.5000 7.8650 2.0100 ;
        RECT  6.4250 0.6800 6.6650 0.8500 ;
        RECT  4.6450 0.6800 4.8850 0.8500 ;
        RECT  3.9250 0.7300 4.0450 1.6200 ;
        RECT  3.7850 1.2300 4.0450 1.3800 ;
        RECT  2.7950 0.6800 3.0350 0.8500 ;
        RECT  1.5150 0.6800 1.7550 0.8000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 11.0200 0.1800 ;
        RECT  9.9650 -0.1800 10.0850 0.6700 ;
        RECT  8.6250 0.4900 8.8650 0.6100 ;
        RECT  8.6250 -0.1800 8.7450 0.6100 ;
        RECT  7.2650 0.4900 7.5050 0.6100 ;
        RECT  7.2650 -0.1800 7.3850 0.6100 ;
        RECT  5.3850 0.4900 5.6250 0.6100 ;
        RECT  5.3850 -0.1800 5.5050 0.6100 ;
        RECT  3.9050 0.4900 4.1450 0.6100 ;
        RECT  3.9050 -0.1800 4.0250 0.6100 ;
        RECT  2.1550 0.4900 2.3950 0.6100 ;
        RECT  2.1550 -0.1800 2.2750 0.6100 ;
        RECT  0.9350 -0.1800 1.0550 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 11.0200 2.7900 ;
        RECT  3.5150 1.9800 3.7550 2.1500 ;
        RECT  3.5150 1.9800 3.6350 2.7900 ;
        RECT  2.6750 1.9800 2.9150 2.1500 ;
        RECT  2.6750 1.9800 2.7950 2.7900 ;
        RECT  1.8350 1.9800 2.0750 2.1500 ;
        RECT  1.8350 1.9800 1.9550 2.7900 ;
        RECT  0.9950 1.9800 1.2350 2.1500 ;
        RECT  0.9950 1.9800 1.1150 2.7900 ;
        RECT  0.2150 1.5600 0.3350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  10.8050 2.2500 4.0250 2.2500 4.0250 2.1500 3.9050 2.1500 3.9050 1.9800 4.1450 1.9800
                 4.1450 2.1300 4.7450 2.1300 4.7450 1.9800 4.9850 1.9800 4.9850 2.1300 5.5850 2.1300
                 5.5850 1.9800 5.8250 1.9800 5.8250 2.1300 6.4250 2.1300 6.4250 1.9800 6.6650 1.9800
                 6.6650 2.1300 7.3250 2.1300 7.3250 1.7400 7.4450 1.7400 7.4450 2.1300 8.1650 2.1300
                 8.1650 1.7400 8.2850 1.7400 8.2850 2.1300 9.0050 2.1300 9.0050 1.7400 9.1250 1.7400
                 9.1250 2.1300 9.8450 2.1300 9.8450 1.7400 9.9650 1.7400 9.9650 2.1300 10.6850 2.1300
                 10.6850 1.5600 10.8050 1.5600 ;
        POLYGON  7.0250 2.0100 6.9050 2.0100 6.9050 1.8600 6.1850 1.8600 6.1850 2.0100 6.0650 2.0100
                 6.0650 1.8600 5.3450 1.8600 5.3450 2.0100 5.2250 2.0100 5.2250 1.8600 4.5050 1.8600
                 4.5050 2.0100 4.3850 2.0100 4.3850 1.8600 3.2750 1.8600 3.2750 2.2100 3.1550 2.2100
                 3.1550 1.8600 2.4350 1.8600 2.4350 2.2100 2.3150 2.2100 2.3150 1.8600 1.5950 1.8600
                 1.5950 2.2100 1.4750 2.2100 1.4750 1.8600 0.7550 1.8600 0.7550 2.2100 0.6350 2.2100
                 0.6350 1.5600 0.7550 1.5600 0.7550 1.7400 1.4750 1.7400 1.4750 1.5600 1.5950 1.5600
                 1.5950 1.7400 2.3150 1.7400 2.3150 1.5600 2.4350 1.5600 2.4350 1.7400 3.1550 1.7400
                 3.1550 1.5600 3.2750 1.5600 3.2750 1.7400 7.0250 1.7400 ;
    END
END AOI222X4

MACRO AOI222X2
    CLASS CORE ;
    FOREIGN AOI222X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9800 0.9900 5.5100 1.1100 ;
        RECT  4.0750 0.9400 5.1000 0.9900 ;
        RECT  4.1300 0.8700 5.1000 0.9900 ;
        RECT  4.0100 0.9900 4.3350 1.0900 ;
        RECT  4.0100 0.9900 4.2500 1.1100 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5300 0.9900 3.8300 1.1100 ;
        RECT  2.9150 0.9400 3.1750 1.1100 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5000 0.9900 1.9600 1.1100 ;
        RECT  0.5950 0.9400 1.6200 1.0300 ;
        RECT  0.7350 0.9100 1.6200 1.0300 ;
        RECT  0.5600 0.9900 0.8550 1.1100 ;
        END
    END A0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7100 1.1100 4.8600 1.5800 ;
        RECT  4.7100 1.1100 4.8300 1.6100 ;
        END
    END C1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2600 1.1500 1.3800 1.6500 ;
        RECT  1.2300 1.1500 1.3800 1.6200 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.2300 3.0900 1.4100 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.8288  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.2700 1.5600 5.3900 2.0100 ;
        RECT  4.4300 1.7300 5.3900 1.8500 ;
        RECT  1.2400 0.6300 4.7300 0.7500 ;
        RECT  4.4300 1.5300 4.5500 2.0100 ;
        RECT  2.2900 1.5300 4.5500 1.6500 ;
        RECT  2.2900 0.6300 2.4100 1.6500 ;
        RECT  2.1000 1.1750 2.4100 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.1900 -0.1800 5.3100 0.6400 ;
        RECT  3.7900 0.3900 4.0300 0.5100 ;
        RECT  3.7900 -0.1800 3.9100 0.5100 ;
        RECT  2.2100 0.3900 2.4500 0.5100 ;
        RECT  2.2100 -0.1800 2.3300 0.5100 ;
        RECT  0.6600 -0.1800 0.7800 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  1.8800 2.0100 2.1200 2.1500 ;
        RECT  1.8800 2.0100 2.0000 2.7900 ;
        RECT  1.0400 2.0100 1.2800 2.1500 ;
        RECT  1.0400 2.0100 1.1600 2.7900 ;
        RECT  0.2600 1.5600 0.3800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.8100 2.2500 2.3900 2.2500 2.3900 2.1500 2.2700 2.1500 2.2700 2.0100 2.5100 2.0100
                 2.5100 2.1300 3.1100 2.1300 3.1100 2.0100 3.3500 2.0100 3.3500 2.1300 4.0100 2.1300
                 4.0100 1.7700 4.1300 1.7700 4.1300 2.1300 4.8500 2.1300 4.8500 1.9700 4.9700 1.9700
                 4.9700 2.1300 5.6900 2.1300 5.6900 1.5600 5.8100 1.5600 ;
        POLYGON  3.7100 2.0100 3.5900 2.0100 3.5900 1.8900 2.8700 1.8900 2.8700 2.0100 2.7500 2.0100
                 2.7500 1.8900 1.6400 1.8900 1.6400 2.2100 1.5200 2.2100 1.5200 1.8900 0.8000 1.8900
                 0.8000 2.2100 0.6800 2.2100 0.6800 1.5600 0.8000 1.5600 0.8000 1.7700 1.5200 1.7700
                 1.5200 1.5600 1.6400 1.5600 1.6400 1.7700 3.7100 1.7700 ;
    END
END AOI222X2

MACRO AOI222X1
    CLASS CORE ;
    FOREIGN AOI222X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9150 1.1750 1.1200 1.4500 ;
        RECT  0.8500 1.2050 1.0350 1.4600 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3000 1.0000 2.5400 1.4400 ;
        RECT  2.3000 1.0000 2.4200 1.4600 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9400 1.2000 2.1800 1.4400 ;
        RECT  1.8100 1.1750 2.0700 1.4350 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.8850 0.5100 1.4400 ;
        RECT  0.3600 0.8850 0.5100 1.3550 ;
        END
    END A0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7150 1.0000 2.8600 1.3450 ;
        RECT  2.6600 1.0850 2.8350 1.4350 ;
        END
    END C1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5550 1.0000 1.6800 1.4600 ;
        RECT  1.5200 1.0000 1.6800 1.4350 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6337  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9700 1.4650 3.1200 1.7250 ;
        RECT  2.9800 0.6500 3.1000 1.7250 ;
        RECT  1.4000 0.7600 3.1000 0.8800 ;
        RECT  2.7200 0.6500 3.1000 0.8800 ;
        RECT  2.6600 1.5600 3.1200 1.6800 ;
        RECT  2.6600 1.5600 2.7800 2.0100 ;
        RECT  1.4000 0.5900 1.5200 0.8800 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.1400 -0.1800 2.2600 0.6400 ;
        RECT  0.3700 -0.1800 0.4900 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  1.0100 1.8200 1.1300 2.7900 ;
        RECT  0.1700 1.5600 0.2900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.2600 2.1500 3.1400 2.1500 3.1400 2.2500 1.4000 2.2500 1.4000 1.8200 1.5200 1.8200
                 1.5200 2.1300 2.2400 2.1300 2.2400 1.5800 2.3600 1.5800 2.3600 2.1300 3.0200 2.1300
                 3.0200 1.8450 3.2600 1.8450 ;
        POLYGON  1.9400 2.0100 1.8200 2.0100 1.8200 1.7000 0.7100 1.7000 0.7100 2.2100 0.5900 2.2100
                 0.5900 1.5600 0.7100 1.5600 0.7100 1.5800 1.8200 1.5800 1.8200 1.5600 1.9400 1.5600 ;
    END
END AOI222X1

MACRO AOI221XL
    CLASS CORE ;
    FOREIGN AOI221XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7350 0.7450 0.9750 0.9350 ;
        RECT  0.5950 0.6500 0.8550 0.8650 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2050 1.0800 2.3250 1.3950 ;
        RECT  2.0450 1.2300 2.3050 1.4200 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.1100 0.5650 1.3800 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 0.9400 2.0150 1.1100 ;
        RECT  1.8050 0.9400 1.9250 1.3250 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 0.9750 1.6350 1.1200 ;
        RECT  1.1750 0.9400 1.4350 1.1200 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3288  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5650 1.1750 2.8300 1.4350 ;
        RECT  2.5650 0.7000 2.6850 1.6600 ;
        RECT  1.3050 0.7000 2.6850 0.8200 ;
        RECT  2.3650 0.4000 2.4850 0.8200 ;
        RECT  1.3050 0.4000 1.4250 0.8200 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.8850 0.4600 2.1250 0.5800 ;
        RECT  1.8850 -0.1800 2.0050 0.5800 ;
        RECT  0.3150 -0.1800 0.4350 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.0150 1.9300 1.1350 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2650 1.9250 1.3250 1.9250 1.3250 1.6000 1.2050 1.6000 1.2050 1.4800 1.4450 1.4800
                 1.4450 1.8050 2.1450 1.8050 2.1450 1.5400 2.2650 1.5400 ;
        POLYGON  1.8450 1.6850 1.7250 1.6850 1.7250 1.5650 1.5650 1.5650 1.5650 1.3600 0.8050 1.3600
                 0.8050 1.6200 0.6550 1.6200 0.6550 1.8300 0.5350 1.8300 0.5350 1.5000 0.6850 1.5000
                 0.6850 1.2400 1.6850 1.2400 1.6850 1.4450 1.8450 1.4450 ;
    END
END AOI221XL

MACRO AOI221X4
    CLASS CORE ;
    FOREIGN AOI221X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 9.2800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6950 0.9900 8.4950 1.1100 ;
        RECT  7.6950 0.9400 7.8150 1.1800 ;
        RECT  7.5550 0.9400 7.8150 1.0900 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1550 0.9900 7.1350 1.1100 ;
        RECT  6.6850 1.2300 6.9450 1.3800 ;
        RECT  6.6850 0.9900 6.8050 1.3800 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5050 0.9900 3.5050 1.1100 ;
        RECT  0.8850 0.9400 1.1450 1.1100 ;
        END
    END A0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9950 1.2300 6.3950 1.3500 ;
        RECT  5.8150 1.2300 6.0750 1.3800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3450 1.2300 2.8650 1.3500 ;
        RECT  1.4650 1.2300 1.7250 1.3800 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2416  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.5750 1.3200 8.6950 2.0100 ;
        RECT  7.7350 1.3200 8.6950 1.4400 ;
        RECT  8.2150 0.6500 8.4550 0.7700 ;
        RECT  1.6250 0.7000 8.3350 0.8200 ;
        RECT  7.7350 1.3200 7.8550 2.0100 ;
        RECT  3.9150 1.5000 7.8550 1.6200 ;
        RECT  7.3750 0.6500 7.6150 0.8200 ;
        RECT  6.3150 0.6500 6.5550 0.8200 ;
        RECT  4.7350 0.6500 4.9750 0.8200 ;
        RECT  3.7850 1.2300 4.0450 1.3800 ;
        RECT  3.9150 0.7000 4.0350 1.6200 ;
        RECT  2.7850 0.6500 3.0250 0.8200 ;
        RECT  1.5050 0.6500 1.7450 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 9.2800 0.1800 ;
        RECT  8.6950 -0.1800 8.8150 0.6400 ;
        RECT  7.7950 0.4600 8.0350 0.5800 ;
        RECT  7.7950 -0.1800 7.9150 0.5800 ;
        RECT  6.9550 0.4600 7.1950 0.5800 ;
        RECT  6.9550 -0.1800 7.0750 0.5800 ;
        RECT  5.4750 0.4600 5.7150 0.5800 ;
        RECT  5.4750 -0.1800 5.5950 0.5800 ;
        RECT  3.8950 0.4600 4.1350 0.5800 ;
        RECT  3.8950 -0.1800 4.0150 0.5800 ;
        RECT  2.1450 0.4600 2.3850 0.5800 ;
        RECT  2.1450 -0.1800 2.2650 0.5800 ;
        RECT  0.9250 -0.1800 1.0450 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 9.2800 2.7900 ;
        RECT  3.5050 1.9800 3.7450 2.1500 ;
        RECT  3.5050 1.9800 3.6250 2.7900 ;
        RECT  2.6650 1.9800 2.9050 2.1500 ;
        RECT  2.6650 1.9800 2.7850 2.7900 ;
        RECT  1.8250 1.9800 2.0650 2.1500 ;
        RECT  1.8250 1.9800 1.9450 2.7900 ;
        RECT  0.9850 1.9800 1.2250 2.1500 ;
        RECT  0.9850 1.9800 1.1050 2.7900 ;
        RECT  0.2050 1.5600 0.3250 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.1150 2.2500 4.0150 2.2500 4.0150 2.1500 3.8950 2.1500 3.8950 1.9800 4.1350 1.9800
                 4.1350 2.1300 4.7350 2.1300 4.7350 1.9800 4.9750 1.9800 4.9750 2.1300 5.5750 2.1300
                 5.5750 1.9800 5.8150 1.9800 5.8150 2.1300 6.4150 2.1300 6.4150 1.9800 6.6550 1.9800
                 6.6550 2.1300 7.3150 2.1300 7.3150 1.7400 7.4350 1.7400 7.4350 2.1300 8.1550 2.1300
                 8.1550 1.5600 8.2750 1.5600 8.2750 2.1300 8.9950 2.1300 8.9950 1.5600 9.1150 1.5600 ;
        POLYGON  7.0150 2.0100 6.8950 2.0100 6.8950 1.8600 6.1750 1.8600 6.1750 2.0100 6.0550 2.0100
                 6.0550 1.8600 5.3350 1.8600 5.3350 2.0100 5.2150 2.0100 5.2150 1.8600 4.4950 1.8600
                 4.4950 2.0100 4.3750 2.0100 4.3750 1.8600 3.2650 1.8600 3.2650 2.2100 3.1450 2.2100
                 3.1450 1.8600 2.4250 1.8600 2.4250 2.2100 2.3050 2.2100 2.3050 1.8600 1.5850 1.8600
                 1.5850 2.2100 1.4650 2.2100 1.4650 1.8600 0.7450 1.8600 0.7450 2.2100 0.6250 2.2100
                 0.6250 1.5600 0.7450 1.5600 0.7450 1.7400 1.4650 1.7400 1.4650 1.5600 1.5850 1.5600
                 1.5850 1.7400 2.3050 1.7400 2.3050 1.5600 2.4250 1.5600 2.4250 1.7400 3.1450 1.7400
                 3.1450 1.5600 3.2650 1.5600 3.2650 1.7400 7.0150 1.7400 ;
    END
END AOI221X4

MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3650 0.9400 4.6250 1.1550 ;
        RECT  4.2450 1.0350 4.4850 1.2250 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3700 0.9900 3.7900 1.1100 ;
        RECT  2.9150 0.9400 3.1750 1.1100 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5000 0.9900 1.9200 1.1100 ;
        RECT  0.5950 0.9400 1.6200 1.0500 ;
        RECT  0.7350 0.9300 1.6200 1.0500 ;
        RECT  0.5200 0.9900 0.8550 1.1100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.1700 1.3800 1.6400 ;
        RECT  1.2400 1.1700 1.3600 1.6700 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 1.2300 3.0500 1.4100 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6208  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3900 1.5300 4.5100 2.0100 ;
        RECT  2.1300 1.5300 4.5100 1.6500 ;
        RECT  4.0300 0.6500 4.2700 0.7700 ;
        RECT  1.3200 0.6900 4.1500 0.8100 ;
        RECT  2.8500 0.6500 3.0900 0.8100 ;
        RECT  2.1300 0.6900 2.2500 1.6500 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.2000 0.6500 1.4400 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  4.5100 -0.1800 4.6300 0.6400 ;
        RECT  3.5500 0.4500 3.7900 0.5700 ;
        RECT  3.5500 -0.1800 3.6700 0.5700 ;
        RECT  2.1500 0.4500 2.3900 0.5700 ;
        RECT  2.1500 -0.1800 2.2700 0.5700 ;
        RECT  0.6200 -0.1800 0.7400 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  1.8400 2.0300 2.0800 2.1500 ;
        RECT  1.8400 2.0300 1.9600 2.7900 ;
        RECT  1.0000 2.0300 1.2400 2.1500 ;
        RECT  1.0000 2.0300 1.1200 2.7900 ;
        RECT  0.2200 1.5600 0.3400 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.9300 2.2500 2.3500 2.2500 2.3500 2.1500 2.2300 2.1500 2.2300 2.0300 2.4700 2.0300
                 2.4700 2.1300 3.0700 2.1300 3.0700 2.0300 3.3100 2.0300 3.3100 2.1300 3.9700 2.1300
                 3.9700 1.7700 4.0900 1.7700 4.0900 2.1300 4.8100 2.1300 4.8100 1.5600 4.9300 1.5600 ;
        POLYGON  3.6700 2.0100 3.5500 2.0100 3.5500 1.9100 2.8300 1.9100 2.8300 2.0100 2.7100 2.0100
                 2.7100 1.9100 1.6000 1.9100 1.6000 2.2100 1.4800 2.2100 1.4800 1.9100 0.7600 1.9100
                 0.7600 2.2100 0.6400 2.2100 0.6400 1.5600 0.7600 1.5600 0.7600 1.7900 1.4800 1.7900
                 1.4800 1.7600 1.6000 1.7600 1.6000 1.7900 2.7100 1.7900 2.7100 1.7700 2.8300 1.7700
                 2.8300 1.7900 3.5500 1.7900 3.5500 1.7700 3.6700 1.7700 ;
    END
END AOI221X2

MACRO AOI221X1
    CLASS CORE ;
    FOREIGN AOI221X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8150 1.0400 1.0900 1.1600 ;
        RECT  0.9400 0.8850 1.0900 1.1600 ;
        RECT  0.8150 1.0400 0.9350 1.2950 ;
        END
    END A1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.2950 2.4800 1.4250 ;
        RECT  2.1000 1.1500 2.2500 1.4350 ;
        END
    END C0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7700 0.5100 1.1450 ;
        RECT  0.3600 0.7700 0.4800 1.3800 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8600 0.9400 1.9800 1.4000 ;
        RECT  1.8100 1.0000 1.9600 1.4350 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 0.9650 1.6700 1.4350 ;
        RECT  1.5400 0.9400 1.6600 1.4400 ;
        END
    END B1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6141  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6400 0.8200 2.7600 2.2050 ;
        RECT  2.4200 0.8200 2.7600 0.9400 ;
        RECT  1.4400 0.7000 2.5600 0.8200 ;
        RECT  2.4400 0.5800 2.5600 0.9400 ;
        RECT  2.3900 0.5950 2.5600 0.8550 ;
        RECT  1.3200 0.6500 1.5600 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.9600 0.4600 2.2000 0.5800 ;
        RECT  1.9600 -0.1800 2.0800 0.5800 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  1.0350 2.1900 1.1550 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.3400 2.2500 1.3800 2.2500 1.3800 1.8000 1.5000 1.8000 1.5000 2.1300 2.2200 2.1300
                 2.2200 1.5550 2.3400 1.5550 ;
        POLYGON  1.9200 2.0100 1.8000 2.0100 1.8000 1.6800 0.6750 1.6800 0.6750 2.2100 0.5550 2.2100
                 0.5550 1.5600 1.8000 1.5600 1.8000 1.5550 1.9200 1.5550 ;
    END
END AOI221X1

MACRO AOI21XL
    CLASS CORE ;
    FOREIGN AOI21XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 0.9800 1.3800 1.4350 ;
        RECT  1.2450 0.9800 1.3650 1.4600 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8250 0.7000 0.9450 1.0200 ;
        RECT  0.6500 0.7000 0.9450 0.9200 ;
        RECT  0.6500 0.5950 0.8000 0.9200 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.9200 0.4750 1.0450 ;
        RECT  0.0700 0.8850 0.2200 1.1500 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1776  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5000 0.8850 1.6700 1.1450 ;
        RECT  1.5000 0.7400 1.6200 1.6750 ;
        RECT  1.4850 1.5550 1.6050 1.7950 ;
        RECT  1.0650 0.7400 1.6200 0.8600 ;
        RECT  1.0650 0.4400 1.1850 0.8600 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  1.4250 0.5000 1.6650 0.6200 ;
        RECT  1.4250 -0.1800 1.5450 0.6200 ;
        RECT  0.3450 -0.1800 0.4650 0.6800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.6150 2.1000 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1850 1.8200 1.0650 1.8200 1.0650 1.7000 0.0750 1.7000 0.0750 1.5800 1.1850 1.5800 ;
    END
END AOI21XL

MACRO AOI21X4
    CLASS CORE ;
    FOREIGN AOI21X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0150 0.9900 4.7550 1.1100 ;
        RECT  4.0750 0.9400 4.3350 1.1100 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 1.1750 3.4100 1.4350 ;
        RECT  3.2550 0.9900 3.3800 1.1800 ;
        RECT  3.2550 0.9400 3.3750 1.1800 ;
        RECT  0.9150 0.9900 3.3800 1.1100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2300 2.7750 1.3500 ;
        RECT  1.1750 1.2300 1.4350 1.3800 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.9664  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.8350 1.3150 4.9550 2.0100 ;
        RECT  4.5950 0.6500 4.8350 0.7700 ;
        RECT  3.7750 1.3150 4.9550 1.4350 ;
        RECT  1.5350 0.7000 4.7150 0.8200 ;
        RECT  3.9950 1.3150 4.1150 2.0100 ;
        RECT  3.7750 1.2300 4.0450 1.4350 ;
        RECT  3.8150 0.5800 3.9350 0.8200 ;
        RECT  3.7750 0.7000 3.8950 1.4350 ;
        RECT  2.6950 0.6500 2.9350 0.8200 ;
        RECT  1.4150 0.6500 1.6550 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  5.0750 -0.1800 5.1950 0.6400 ;
        RECT  4.1750 0.4600 4.4150 0.5800 ;
        RECT  4.1750 -0.1800 4.2950 0.5800 ;
        RECT  3.3350 0.4600 3.5750 0.5800 ;
        RECT  3.3350 -0.1800 3.4550 0.5800 ;
        RECT  2.0550 0.4600 2.2950 0.5800 ;
        RECT  2.0550 -0.1800 2.1750 0.5800 ;
        RECT  0.8350 -0.1800 0.9550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  3.0950 1.7950 3.3350 2.1500 ;
        RECT  3.0950 1.7950 3.2150 2.7900 ;
        RECT  2.2550 1.7950 2.4950 2.1500 ;
        RECT  2.2550 1.7950 2.3750 2.7900 ;
        RECT  1.4150 1.7950 1.6550 2.1500 ;
        RECT  1.4150 1.7950 1.5350 2.7900 ;
        RECT  0.5750 1.7950 0.8150 2.1500 ;
        RECT  0.5750 1.7950 0.6950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.3750 2.2500 3.5750 2.2500 3.5750 1.6750 2.8550 1.6750 2.8550 2.2100 2.7350 2.2100
                 2.7350 1.6750 2.0150 1.6750 2.0150 2.2100 1.8950 2.2100 1.8950 1.6750 1.1750 1.6750
                 1.1750 2.2100 1.0550 2.2100 1.0550 1.6750 0.3350 1.6750 0.3350 2.2100 0.2150 2.2100
                 0.2150 1.5550 3.6950 1.5550 3.6950 2.1300 4.4150 2.1300 4.4150 1.5600 4.5350 1.5600
                 4.5350 2.1300 5.2550 2.1300 5.2550 1.5600 5.3750 1.5600 ;
    END
END AOI21X4

MACRO AOI21X2
    CLASS CORE ;
    FOREIGN AOI21X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4832  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3300 1.2500 2.4500 2.0100 ;
        RECT  2.1300 1.2500 2.4500 1.3700 ;
        RECT  2.1300 0.6200 2.2500 1.3700 ;
        RECT  2.1000 0.7400 2.2500 1.1450 ;
        RECT  1.1300 0.7400 2.2500 0.8600 ;
        RECT  1.0100 0.6900 1.2500 0.8100 ;
        END
    END Y
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.2200 1.2150 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 0.9800 1.6900 1.2200 ;
        RECT  1.5200 0.9800 1.6700 1.4350 ;
        RECT  0.6450 0.9800 1.6900 1.1000 ;
        RECT  0.5100 1.0100 0.7650 1.1300 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.8200 2.8850 1.0900 ;
        RECT  2.3700 0.8800 2.7450 1.1300 ;
        END
    END B0
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  1.4900 1.7950 1.6100 2.7900 ;
        RECT  0.6500 1.7950 0.7700 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.5500 -0.1800 2.6700 0.6800 ;
        RECT  1.6500 0.5000 1.8900 0.6200 ;
        RECT  1.6500 -0.1800 1.7700 0.6200 ;
        RECT  0.4300 -0.1800 0.5500 0.6800 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  2.8700 2.2500 1.9100 2.2500 1.9100 1.6750 1.1900 1.6750 1.1900 2.2100 1.0700 2.2100
                 1.0700 1.6750 0.3500 1.6750 0.3500 2.2100 0.2300 2.2100 0.2300 1.5550 2.0300 1.5550
                 2.0300 2.1300 2.7500 2.1300 2.7500 1.5600 2.8700 1.5600 ;
    END
END AOI21X2

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9700 1.0550 1.2100 1.1950 ;
        RECT  0.9400 1.1500 1.0900 1.4350 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0200 0.8200 1.4350 ;
        RECT  0.7000 1.0050 0.8200 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.8250 0.5100 1.2800 ;
        RECT  0.3800 0.8250 0.5000 1.3050 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3196  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 0.8850 1.6700 1.1450 ;
        RECT  1.3950 0.7650 1.5150 2.2100 ;
        RECT  0.8600 0.7650 1.5150 0.8850 ;
        RECT  0.8600 0.6450 0.9800 0.8850 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  1.2200 0.5250 1.4600 0.6450 ;
        RECT  1.2200 -0.1800 1.3400 0.6450 ;
        RECT  0.2200 -0.1800 0.3400 0.7050 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.5550 1.7950 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.0950 2.2100 0.9750 2.2100 0.9750 1.6750 0.2550 1.6750 0.2550 2.2100 0.1350 2.2100
                 0.1350 1.5550 1.0950 1.5550 ;
    END
END AOI21X1

MACRO AOI211XL
    CLASS CORE ;
    FOREIGN AOI211XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3300 1.0550 1.4750 1.2950 ;
        RECT  1.2300 1.1750 1.4000 1.4350 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8700 1.0550 1.1100 1.2600 ;
        RECT  0.9400 1.0550 1.0900 1.4500 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.1600 0.7500 1.2900 ;
        RECT  0.3600 1.1600 0.5100 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1200 0.8900 0.2400 1.3500 ;
        RECT  0.0700 0.8850 0.2200 1.3200 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2448  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6150 0.5150 1.7350 1.9300 ;
        RECT  1.5200 1.4650 1.7350 1.7250 ;
        RECT  0.7750 0.8150 1.7350 0.9350 ;
        RECT  0.7750 0.5150 0.8950 0.9350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  1.1350 0.5750 1.3750 0.6950 ;
        RECT  1.1350 -0.1800 1.2550 0.6950 ;
        RECT  0.1350 -0.1800 0.2550 0.7550 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  0.5550 1.8100 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1550 1.8700 0.9150 1.8700 0.9150 1.6900 0.3150 1.6900 0.3150 1.8700 0.0750 1.8700
                 0.0750 1.7500 0.1950 1.7500 0.1950 1.5700 1.0350 1.5700 1.0350 1.7500 1.1550 1.7500 ;
    END
END AOI211XL

MACRO AOI211X4
    CLASS CORE ;
    FOREIGN AOI211X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4350 0.9900 3.4350 1.1100 ;
        RECT  0.5950 0.9400 0.8550 1.1100 ;
        END
    END A0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5450 0.9400 6.6650 1.1800 ;
        RECT  5.9650 0.9900 6.6650 1.1100 ;
        RECT  6.3950 0.9400 6.6650 1.1100 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3650 0.9700 5.0250 1.0900 ;
        RECT  4.3650 0.9400 4.6250 1.0900 ;
        RECT  4.2850 0.9900 4.5250 1.1100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2750 1.2300 2.7950 1.3500 ;
        RECT  2.3350 1.2300 2.5950 1.3800 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2416  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.8050 1.3000 6.9250 2.0100 ;
        RECT  5.9650 1.3000 6.9250 1.4200 ;
        RECT  6.5450 0.6500 6.7850 0.7700 ;
        RECT  1.5550 0.7000 6.6650 0.8200 ;
        RECT  5.9650 1.2300 6.0850 2.0100 ;
        RECT  4.0250 1.2300 6.0850 1.3500 ;
        RECT  5.7050 0.6500 5.9450 0.8200 ;
        RECT  4.8650 0.6500 5.1050 0.8200 ;
        RECT  4.0250 0.6500 4.2650 0.8200 ;
        RECT  4.0250 0.6500 4.1450 1.3500 ;
        RECT  3.7850 0.9400 4.1450 1.0900 ;
        RECT  2.7150 0.6500 2.9550 0.8200 ;
        RECT  1.4350 0.6500 1.6750 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  7.0250 -0.1800 7.1450 0.6400 ;
        RECT  6.1250 0.4600 6.3650 0.5800 ;
        RECT  6.1250 -0.1800 6.2450 0.5800 ;
        RECT  5.2850 0.4600 5.5250 0.5800 ;
        RECT  5.2850 -0.1800 5.4050 0.5800 ;
        RECT  4.4450 0.4600 4.6850 0.5800 ;
        RECT  4.4450 -0.1800 4.5650 0.5800 ;
        RECT  3.6050 0.4600 3.8450 0.5800 ;
        RECT  3.6050 -0.1800 3.7250 0.5800 ;
        RECT  2.0750 0.4600 2.3150 0.5800 ;
        RECT  2.0750 -0.1800 2.1950 0.5800 ;
        RECT  0.8550 -0.1800 0.9750 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  3.5550 2.0700 3.6750 2.7900 ;
        RECT  2.6550 1.7400 2.7750 2.7900 ;
        RECT  1.8150 1.7400 1.9350 2.7900 ;
        RECT  0.9750 1.7400 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.3450 2.2500 3.9250 2.2500 3.9250 1.8600 3.8050 1.8600 3.8050 1.7400 4.0450 1.7400
                 4.0450 2.1300 4.7050 2.1300 4.7050 1.7400 4.8250 1.7400 4.8250 2.1300 5.5450 2.1300
                 5.5450 1.4700 5.6650 1.4700 5.6650 2.1300 6.3850 2.1300 6.3850 1.5400 6.5050 1.5400
                 6.5050 2.1300 7.2250 2.1300 7.2250 1.4700 7.3450 1.4700 ;
        POLYGON  5.2450 2.0100 5.1250 2.0100 5.1250 1.6200 4.4050 1.6200 4.4050 2.0100 4.2850 2.0100
                 4.2850 1.6200 3.1950 1.6200 3.1950 2.2100 3.0750 2.2100 3.0750 1.6200 2.3550 1.6200
                 2.3550 2.2100 2.2350 2.2100 2.2350 1.6200 1.5150 1.6200 1.5150 2.2100 1.3950 2.2100
                 1.3950 1.6200 0.6750 1.6200 0.6750 2.2100 0.5550 2.2100 0.5550 1.5000 4.2850 1.5000
                 4.2850 1.4700 4.4050 1.4700 4.4050 1.5000 5.1250 1.5000 5.1250 1.4700 5.2450 1.4700 ;
    END
END AOI211X4

MACRO AOI211X2
    CLASS CORE ;
    FOREIGN AOI211X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.0600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2050 0.9400 3.5250 1.1600 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9400 2.8850 1.1550 ;
        RECT  2.5050 0.9400 2.8850 1.1300 ;
        END
    END B0
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5550 0.9900 1.7950 1.1100 ;
        RECT  0.5950 0.9400 1.6750 1.0600 ;
        RECT  0.4350 0.9900 0.8550 1.1100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0550 1.1800 1.4350 1.4000 ;
        END
    END A1
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6208  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.3850 1.2800 3.5050 1.9900 ;
        RECT  2.2650 1.2800 3.5050 1.4000 ;
        RECT  3.1250 0.6500 3.3650 0.7700 ;
        RECT  1.1950 0.7000 3.2450 0.8200 ;
        RECT  2.2650 0.6500 2.5050 0.8200 ;
        RECT  2.2650 0.6500 2.3850 1.4000 ;
        RECT  2.1000 0.7000 2.3850 1.1450 ;
        RECT  1.0750 0.6500 1.3150 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.0600 0.1800 ;
        RECT  3.6050 -0.1800 3.7250 0.6400 ;
        RECT  2.6850 0.4600 2.9250 0.5800 ;
        RECT  2.6850 -0.1800 2.8050 0.5800 ;
        RECT  1.8450 0.4600 2.0850 0.5800 ;
        RECT  1.8450 -0.1800 1.9650 0.5800 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.0600 2.7900 ;
        RECT  1.8750 2.1400 1.9950 2.7900 ;
        RECT  0.9750 1.7600 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.9250 2.2300 2.1850 2.2300 2.1850 1.8800 2.0650 1.8800 2.0650 1.7600 2.3050 1.7600
                 2.3050 2.1100 2.9650 2.1100 2.9650 1.5200 3.0850 1.5200 3.0850 2.1100 3.8050 2.1100
                 3.8050 1.3400 3.9250 1.3400 ;
        POLYGON  2.6650 1.9900 2.5450 1.9900 2.5450 1.6400 1.5150 1.6400 1.5150 2.2100 1.3950 2.2100
                 1.3950 1.6400 0.6750 1.6400 0.6750 2.2100 0.5550 2.2100 0.5550 1.5200 2.6650 1.5200 ;
    END
END AOI211X2

MACRO AOI211X1
    CLASS CORE ;
    FOREIGN AOI211X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.0950 1.6700 1.4350 ;
        RECT  1.4800 0.9750 1.6000 1.3150 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.0100 1.1800 1.1500 ;
        RECT  0.9400 1.0100 1.0900 1.4350 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.9800 0.8000 1.4350 ;
        RECT  0.6800 0.9600 0.8000 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7800 0.5100 1.1500 ;
        RECT  0.3200 0.8150 0.4400 1.1900 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.4400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6400 1.5550 1.9100 1.6750 ;
        RECT  1.7900 0.7200 1.9100 1.6750 ;
        RECT  0.8600 0.7200 1.9100 0.8400 ;
        RECT  1.6400 1.5550 1.7600 2.2100 ;
        RECT  1.5200 0.6000 1.7600 0.8400 ;
        RECT  1.5200 0.5950 1.6700 0.8550 ;
        RECT  0.7400 0.6700 0.9800 0.7900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  1.1600 0.4800 1.4000 0.6000 ;
        RECT  1.1600 -0.1800 1.2800 0.6000 ;
        RECT  0.1600 -0.1800 0.2800 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  0.5800 1.7950 0.7000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1200 2.2100 1.0000 2.2100 1.0000 1.6750 0.2800 1.6750 0.2800 2.2100 0.1600 2.2100
                 0.1600 1.5550 1.1200 1.5550 ;
    END
END AOI211X1

MACRO AO22XL
    CLASS CORE ;
    FOREIGN AO22XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8850 0.8200 1.3200 ;
        RECT  0.7000 0.8600 0.8200 1.3200 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9800 1.0900 1.1600 1.3300 ;
        RECT  0.9400 1.1750 1.1450 1.4350 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0300 0.5100 1.5000 ;
        RECT  0.3600 1.0300 0.4800 1.5300 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4650 1.9600 1.8100 ;
        RECT  1.5200 1.4650 1.9600 1.5850 ;
        RECT  1.5200 1.4100 1.8000 1.5850 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 1.4000 2.8250 1.5200 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.3900 0.8850 2.5100 1.5200 ;
        RECT  2.1600 0.8850 2.5400 1.0250 ;
        RECT  2.1600 0.6700 2.2800 1.0250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.6800 0.7300 1.9200 0.8500 ;
        RECT  1.6800 -0.1800 1.8000 0.8500 ;
        RECT  0.2000 -0.1800 0.3200 0.9100 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.2050 1.9800 2.3250 2.7900 ;
        RECT  0.5550 1.8900 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.0400 1.3100 1.9200 1.3100 1.9200 1.2900 1.4000 1.2900 1.4000 1.7050 1.5150 1.7050
                 1.5150 2.0100 1.3950 2.0100 1.3950 1.8250 1.2800 1.8250 1.2800 0.9700 1.0600 0.9700
                 1.0600 0.8500 0.9400 0.8500 0.9400 0.7300 1.1800 0.7300 1.1800 0.8500 1.4000 0.8500
                 1.4000 1.1700 1.9200 1.1700 1.9200 1.0700 2.0400 1.0700 ;
        POLYGON  1.9950 2.0700 1.8750 2.0700 1.8750 2.2500 0.9750 2.2500 0.9750 1.7700 0.3150 1.7700
                 0.3150 1.9500 0.0750 1.9500 0.0750 1.8300 0.1950 1.8300 0.1950 1.6500 1.0950 1.6500
                 1.0950 2.1300 1.7550 2.1300 1.7550 1.9500 1.9950 1.9500 ;
    END
END AO22XL

MACRO AO22X4
    CLASS CORE ;
    FOREIGN AO22X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.0600 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 0.8150 0.8200 1.2350 ;
        RECT  0.7000 0.7950 0.8200 1.2350 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0550 0.9050 1.1750 1.2350 ;
        RECT  0.9400 0.8850 1.0900 1.2150 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7600 0.5100 1.2100 ;
        RECT  0.3800 0.7600 0.5000 1.2350 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7550 1.2300 2.0150 1.3800 ;
        RECT  1.5350 1.1700 1.8750 1.2900 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.4050 1.1750 3.7000 1.4350 ;
        RECT  2.5450 1.3200 3.5250 1.4400 ;
        RECT  3.4050 0.6900 3.5250 1.4400 ;
        RECT  3.3850 1.3200 3.5050 2.2100 ;
        RECT  2.1550 0.6900 3.5250 0.8100 ;
        RECT  2.9950 0.6500 3.2350 0.8100 ;
        RECT  2.5450 1.3200 2.6650 2.2100 ;
        RECT  2.0350 0.6500 2.2750 0.7700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.0600 0.1800 ;
        RECT  3.4750 0.4500 3.7150 0.5700 ;
        RECT  3.4750 -0.1800 3.5950 0.5700 ;
        RECT  2.5150 0.4500 2.7550 0.5700 ;
        RECT  2.5150 -0.1800 2.6350 0.5700 ;
        RECT  1.6750 -0.1800 1.7950 0.6400 ;
        RECT  0.2200 -0.1800 0.3400 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.0600 2.7900 ;
        RECT  3.8050 1.5600 3.9250 2.7900 ;
        RECT  2.9650 1.5600 3.0850 2.7900 ;
        RECT  2.0650 2.2300 2.1850 2.7900 ;
        RECT  0.5550 1.5950 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.2850 1.0900 3.0450 1.0900 3.0450 1.0500 2.5350 1.0500 2.5350 1.1100 2.2950 1.1100
                 2.2950 1.0500 1.4150 1.0500 1.4150 1.4100 1.5150 1.4100 1.5150 2.0100 1.3950 2.0100
                 1.3950 1.5300 1.2950 1.5300 1.2950 0.6750 0.9150 0.6750 0.9150 0.5550 1.4150 0.5550
                 1.4150 0.9300 3.1650 0.9300 3.1650 0.9700 3.2850 0.9700 ;
        POLYGON  1.9350 2.2500 0.9750 2.2500 0.9750 1.4750 0.2550 1.4750 0.2550 2.0800 0.1350 2.0800
                 0.1350 1.3550 1.0950 1.3550 1.0950 2.1300 1.8150 2.1300 1.8150 1.5000 1.9350 1.5000 ;
    END
END AO22X4

MACRO AO22X2
    CLASS CORE ;
    FOREIGN AO22X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9350 0.9900 1.0550 1.2300 ;
        RECT  0.6500 0.9900 1.0550 1.1100 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3150 0.8900 1.4350 1.2550 ;
        RECT  1.1750 0.8900 1.4350 1.1000 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.9850 0.4150 1.4400 ;
        RECT  0.2950 0.9650 0.4150 1.4400 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7950 1.0200 1.9600 1.4400 ;
        RECT  1.7950 1.0000 1.9150 1.4400 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6650 1.1450 2.7850 2.2100 ;
        RECT  2.4200 1.1450 2.7850 1.2650 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.3750 0.5900 2.4950 1.0250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  2.7950 -0.1800 2.9150 0.6400 ;
        RECT  1.9550 -0.1800 2.0750 0.6400 ;
        RECT  0.4100 -0.1800 0.5300 0.8300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  3.0850 1.5600 3.2050 2.7900 ;
        RECT  2.1850 2.0100 2.4250 2.1500 ;
        RECT  2.1850 2.0100 2.3050 2.7900 ;
        RECT  0.6150 2.0800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2550 1.1500 2.1350 1.1500 2.1350 0.8800 1.6750 0.8800 1.6750 1.5600 1.6950 1.5600
                 1.6950 1.6800 1.4550 1.6800 1.4550 1.5600 1.5550 1.5600 1.5550 0.7700 1.0350 0.7700
                 1.0350 0.6500 1.6750 0.6500 1.6750 0.7600 2.2550 0.7600 ;
        POLYGON  2.0550 1.9200 1.0950 1.9200 1.0950 1.6800 0.0750 1.6800 0.0750 1.5600 1.2150 1.5600
                 1.2150 1.8000 1.9350 1.8000 1.9350 1.5600 2.0550 1.5600 ;
    END
END AO22X2

MACRO AO22X1
    CLASS CORE ;
    FOREIGN AO22X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9350 0.9100 1.0550 1.1500 ;
        RECT  0.6500 0.9100 1.0550 1.0300 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 0.9400 1.4350 1.1500 ;
        RECT  1.2750 0.9400 1.3950 1.3050 ;
        END
    END B1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.0300 0.4150 1.3700 ;
        RECT  0.2950 0.9500 0.4150 1.3700 ;
        RECT  0.0700 1.0300 0.2200 1.4400 ;
        END
    END A0
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.7950 1.0150 1.9600 1.4350 ;
        RECT  1.7950 1.0000 1.9150 1.4400 ;
        END
    END B0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6450 1.1450 2.7650 2.2100 ;
        RECT  2.4200 1.1450 2.7650 1.2650 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  2.3750 0.5900 2.4950 1.0250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.9550 -0.1800 2.0750 0.6400 ;
        RECT  0.4100 -0.1800 0.5300 0.8300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.1650 2.0100 2.4050 2.1500 ;
        RECT  2.1650 2.0100 2.2850 2.7900 ;
        RECT  0.6150 2.0800 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2550 1.1500 2.1350 1.1500 2.1350 0.8800 1.6750 0.8800 1.6750 1.6200 1.4350 1.6200
                 1.4350 1.5000 1.5550 1.5000 1.5550 0.7700 1.0150 0.7700 1.0150 0.6500 1.6750 0.6500
                 1.6750 0.7600 2.2550 0.7600 ;
        POLYGON  2.0350 1.8600 1.0750 1.8600 1.0750 1.6800 0.0750 1.6800 0.0750 1.5600 1.1950 1.5600
                 1.1950 1.7400 1.9150 1.7400 1.9150 1.5600 2.0350 1.5600 ;
    END
END AO22X1

MACRO AO21XL
    CLASS CORE ;
    FOREIGN AO21XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.4000 1.6700 1.7350 ;
        RECT  1.4000 1.3550 1.6400 1.5200 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.2000 1.1700 1.3200 ;
        RECT  1.0500 1.0800 1.1700 1.3200 ;
        RECT  0.6500 1.1750 0.8000 1.4350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0650 0.5300 1.5000 ;
        RECT  0.4100 1.0400 0.5300 1.5000 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1300 1.4000 2.8250 1.5200 ;
        RECT  2.1300 0.6800 2.2500 1.5200 ;
        RECT  2.1000 0.8850 2.2500 1.1450 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  1.6500 0.7400 1.8900 0.8600 ;
        RECT  1.6500 -0.1800 1.7700 0.8600 ;
        RECT  0.5500 -0.1800 0.6700 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.1800 1.9800 2.3000 2.7900 ;
        RECT  0.8000 1.8600 0.9200 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9700 1.2400 1.9100 1.2400 1.9100 1.9800 1.7900 1.9800 1.7900 1.1000 1.2900 1.1000
                 1.2900 0.6800 1.4100 0.6800 1.4100 0.9800 1.9100 0.9800 1.9100 1.0000 1.9700 1.0000 ;
        POLYGON  1.4000 1.9200 1.1600 1.9200 1.1600 1.7400 0.5600 1.7400 0.5600 1.9200 0.3200 1.9200
                 0.3200 1.8000 0.4400 1.8000 0.4400 1.6200 1.2800 1.6200 1.2800 1.8000 1.4000 1.8000 ;
    END
END AO21XL

MACRO AO21X4
    CLASS CORE ;
    FOREIGN AO21X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.0700 1.1550 1.4350 ;
        RECT  1.0350 1.0650 1.1550 1.4350 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0250 0.8200 1.4600 ;
        RECT  0.7000 1.0000 0.8200 1.4600 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 0.7600 0.5100 1.2250 ;
        RECT  0.3800 0.7600 0.5000 1.2500 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2600 0.8850 3.4100 1.1450 ;
        RECT  2.9800 0.8850 3.4100 1.0050 ;
        RECT  2.9800 0.7600 3.1000 1.6800 ;
        RECT  2.9650 1.5600 3.0850 2.2100 ;
        RECT  2.1250 1.3200 3.1000 1.4400 ;
        RECT  1.8800 0.7600 3.1000 0.8800 ;
        RECT  2.5400 0.5900 2.6600 0.8800 ;
        RECT  2.1250 1.3200 2.2450 2.2100 ;
        RECT  1.7000 0.7100 2.0000 0.8300 ;
        RECT  1.7000 0.5900 1.8200 0.8300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  2.9600 -0.1800 3.0800 0.6400 ;
        RECT  2.1200 -0.1800 2.2400 0.6400 ;
        RECT  1.2800 -0.1800 1.4000 0.6400 ;
        RECT  0.2200 -0.1800 0.3400 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.3850 1.5600 3.5050 2.7900 ;
        RECT  2.5450 1.5600 2.6650 2.7900 ;
        RECT  1.7050 1.9700 1.8250 2.7900 ;
        RECT  0.4950 1.8200 0.7350 2.1450 ;
        RECT  0.4950 1.8200 0.6150 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.8600 1.1900 1.5150 1.1900 1.5150 1.8200 1.3950 1.8200 1.3950 0.8800 0.8600 0.8800
                 0.8600 0.5900 0.9800 0.5900 0.9800 0.7600 1.5150 0.7600 1.5150 1.0700 2.8600 1.0700 ;
        POLYGON  1.0950 2.2050 0.9750 2.2050 0.9750 1.7000 0.2550 1.7000 0.2550 2.2050 0.1350 2.2050
                 0.1350 1.5550 0.2550 1.5550 0.2550 1.5800 0.9750 1.5800 0.9750 1.5550 1.0950 1.5550 ;
    END
END AO21X4

MACRO AO21X2
    CLASS CORE ;
    FOREIGN AO21X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2250 1.0000 1.3800 1.4600 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8350 0.9900 0.9550 1.2300 ;
        RECT  0.6500 0.9900 0.9550 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0650 0.5100 1.5200 ;
        RECT  0.3900 0.9500 0.5100 1.5200 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2250 1.2950 2.3450 2.2100 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  1.9750 1.0550 2.2200 1.1750 ;
        RECT  1.9750 0.5900 2.0950 1.1750 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  2.3950 -0.1800 2.5150 0.6400 ;
        RECT  1.5550 -0.1800 1.6750 0.6400 ;
        RECT  0.3350 -0.1800 0.4550 0.8300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.6450 1.5600 2.7650 2.7900 ;
        RECT  1.8050 1.9700 1.9250 2.7900 ;
        RECT  0.6150 2.1000 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.8550 1.2300 1.6200 1.2300 1.6200 1.7000 1.6150 1.7000 1.6150 1.8200 1.4950 1.8200
                 1.4950 1.5800 1.5000 1.5800 1.5000 0.8800 1.0750 0.8800 1.0750 0.5900 1.1950 0.5900
                 1.1950 0.7600 1.6200 0.7600 1.6200 0.9900 1.8550 0.9900 ;
        RECT  0.0750 1.6400 1.2550 1.7600 ;
    END
END AO21X2

MACRO AO21X1
    CLASS CORE ;
    FOREIGN AO21X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2050 1.1050 1.3800 1.4350 ;
        RECT  1.1950 1.0000 1.3400 1.3250 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 0.7200 0.8800 0.9600 ;
        RECT  0.6500 0.5950 0.8400 0.8550 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.7600 0.5100 1.2600 ;
        RECT  0.3600 0.7600 0.5100 1.2300 ;
        END
    END A0
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1500 1.2950 2.2700 2.2100 ;
        RECT  1.8100 1.2950 2.2700 1.4150 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        RECT  1.8400 0.5900 1.9600 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.4200 -0.1800 1.5400 0.6400 ;
        RECT  0.2600 -0.1800 0.3800 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.7300 1.9450 1.8500 2.7900 ;
        RECT  0.5800 1.6200 0.7000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6800 1.2300 1.6200 1.2300 1.6200 1.6750 1.5400 1.6750 1.5400 1.7950 1.4200 1.7950
                 1.4200 1.5550 1.5000 1.5550 1.5000 0.8800 1.0000 0.8800 1.0000 0.4000 1.1200 0.4000
                 1.1200 0.7600 1.6200 0.7600 1.6200 0.9900 1.6800 0.9900 ;
        POLYGON  1.1800 1.6800 0.8200 1.6800 0.8200 1.5000 0.3400 1.5000 0.3400 1.6800 0.1000 1.6800
                 0.1000 1.5600 0.2200 1.5600 0.2200 1.3800 0.9400 1.3800 0.9400 1.5600 1.1800 1.5600 ;
    END
END AO21X1

MACRO ANTENNA
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN ANTENNA 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116 LAYER Metal1 ;
#   ANTENNAGATEAREA 0.00001  LAYER Metal1  ;
    
    PORT
      LAYER Metal1 ;
	RECT 0.185 0.3 0.685 2.31 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
	RECT 0 -0.18 0.87 0.18 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
	RECT 0 2.43 0.87 2.79 ;
    END
  END VDD
END ANTENNA


#MACRO ANTENNA
#    CLASS CORE ;
#    FOREIGN ANTENNA 0 0 ;
#   ORIGIN 0.0000 0.0000 ;
#    SIZE 0.8700 BY 2.6100 ;
#    SYMMETRY X Y ;
#   SITE gsclib090site ;
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNADIFFAREA 1.1160  LAYER Metal1  ;
#        ANTENNAGATEAREA 0.00001  LAYER Metal1  ;
#        PORT
#        LAYER Metal1 ;
#        RECT  0.1850 0.3000 0.6850 2.3100 ;
#        END
#    END A
#    PIN VSS
#	 DIRECTION INPUT ;
#	 USE ground ;
#	 SHAPE ABUTMENT ;
#	 PORT
#	 LAYER Metal1 ;
#	 RECT  0.0000 -0.1800 0.8700 0.1800 ;
#	 END
#    END VSS
#    PIN VDD
#	 DIRECTION INPUT ;
#	 USE power ;
#	 SHAPE ABUTMENT ;
#	 PORT
#	 LAYER Metal1 ;
#        RECT  0.0000 2.4300 0.8700 2.7900 ;
#        END
#    END VDD
#END ANTENNA

MACRO AND4XL
    CLASS CORE ;
    FOREIGN AND4XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.2300 0.5650 1.5000 ;
        RECT  0.3250 1.1000 0.5650 1.5000 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8150 1.0950 1.0900 1.4600 ;
        RECT  0.8150 1.0950 0.9350 1.4650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2100 1.0950 1.3800 1.5600 ;
        RECT  1.2100 1.0950 1.3300 1.5900 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.3700 1.9600 1.7250 ;
        RECT  1.7400 1.2150 1.8600 1.5750 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3550 0.8550 2.4750 1.8300 ;
        RECT  2.1300 0.8550 2.4750 0.9750 ;
        RECT  2.1000 0.5950 2.2500 0.8550 ;
        RECT  1.9350 0.5950 2.2500 0.7350 ;
        RECT  1.9350 0.4950 2.0550 0.7350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.5150 -0.1800 1.6350 0.7350 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.8750 2.2300 1.9950 2.7900 ;
        RECT  0.9150 2.2300 1.0350 2.7900 ;
        RECT  0.1350 1.7100 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.9800 1.0950 1.8600 1.0950 1.8600 0.9750 1.6200 0.9750 1.6200 1.8300 1.5150 1.8300
                 1.5150 1.9500 1.3950 1.9500 1.3950 1.8300 0.4950 1.8300 0.4950 1.7100 1.5000 1.7100
                 1.5000 0.9750 0.3950 0.9750 0.3950 0.6750 0.2750 0.6750 0.2750 0.5550 0.5150 0.5550
                 0.5150 0.8550 1.9800 0.8550 ;
    END
END AND4XL

MACRO AND4X8
    CLASS CORE ;
    FOREIGN AND4X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.2500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8400 0.9700 2.0800 1.0900 ;
        RECT  1.8400 0.5950 1.9600 1.0900 ;
        RECT  1.8100 0.5950 1.9600 0.8550 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9400 2.8850 1.0900 ;
        RECT  1.2950 1.2100 2.7800 1.3300 ;
        RECT  2.6600 0.9400 2.7800 1.3300 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0200 1.1050 3.2950 1.3450 ;
        RECT  0.9400 1.4500 3.1400 1.5700 ;
        RECT  3.0200 1.1050 3.1400 1.5700 ;
        RECT  0.9400 1.1750 1.0900 1.5700 ;
        RECT  0.7550 1.2800 1.0900 1.4000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.4950 1.6900 3.6150 1.8100 ;
        RECT  3.4950 1.2200 3.6150 1.8100 ;
        RECT  3.2600 1.4650 3.6150 1.8100 ;
        RECT  0.4950 1.2200 0.6150 1.8100 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9150 1.2750 7.0350 2.2100 ;
        RECT  4.3950 1.2750 7.0350 1.3950 ;
        RECT  6.5950 0.7150 6.8350 0.8350 ;
        RECT  4.1350 0.7650 6.7150 0.8850 ;
        RECT  6.0750 1.1750 6.3100 1.4350 ;
        RECT  6.0750 0.7650 6.1950 2.2100 ;
        RECT  5.7550 0.7150 5.9950 0.8850 ;
        RECT  5.2350 1.2750 5.3550 2.2100 ;
        RECT  4.9150 0.7150 5.1550 0.8850 ;
        RECT  4.3950 1.2750 4.5150 2.2100 ;
        RECT  4.0150 0.7150 4.2550 0.8350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.2500 0.1800 ;
        RECT  6.2350 -0.1800 6.3550 0.6450 ;
        RECT  5.3950 -0.1800 5.5150 0.6450 ;
        RECT  4.4950 -0.1800 4.6150 0.6400 ;
        RECT  3.5950 0.4600 3.8350 0.5800 ;
        RECT  3.5950 -0.1800 3.7150 0.5800 ;
        RECT  0.3350 -0.1800 0.4550 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.2500 2.7900 ;
        RECT  6.4950 1.5150 6.6150 2.7900 ;
        RECT  5.6550 1.5150 5.7750 2.7900 ;
        RECT  4.8150 1.5150 4.9350 2.7900 ;
        RECT  3.8550 2.1700 4.0950 2.2900 ;
        RECT  3.8550 2.1700 3.9750 2.7900 ;
        RECT  2.8950 2.1700 3.1350 2.2900 ;
        RECT  2.8950 2.1700 3.0150 2.7900 ;
        RECT  1.9350 2.1700 2.1750 2.2900 ;
        RECT  1.9350 2.1700 2.0550 2.7900 ;
        RECT  0.9750 2.1700 1.2150 2.2900 ;
        RECT  0.9750 2.1700 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.7150 1.1550 3.8550 1.1550 3.8550 2.0500 3.5550 2.0500 3.5550 2.2100 3.4350 2.2100
                 3.4350 2.0500 2.5950 2.0500 2.5950 2.2100 2.4750 2.2100 2.4750 2.0500 1.6350 2.0500
                 1.6350 2.2100 1.5150 2.2100 1.5150 2.0500 0.6750 2.0500 0.6750 2.2100 0.5550 2.2100
                 0.5550 1.9300 3.7350 1.9300 3.7350 0.8200 2.2400 0.8200 2.2400 0.7700 2.1200 0.7700
                 2.1200 0.6500 2.3600 0.6500 2.3600 0.7000 3.8550 0.7000 3.8550 1.0350 5.7150 1.0350 ;
    END
END AND4X8

MACRO AND4X6
    CLASS CORE ;
    FOREIGN AND4X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.3800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8400 0.9700 2.0800 1.0900 ;
        RECT  1.8400 0.5950 1.9600 1.0900 ;
        RECT  1.8100 0.5950 1.9600 0.8550 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.6250 0.9400 2.8850 1.0900 ;
        RECT  1.3000 1.2100 2.7800 1.3300 ;
        RECT  2.6600 0.9400 2.7800 1.3300 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.4500 3.3000 1.5700 ;
        RECT  3.1800 1.2200 3.3000 1.5700 ;
        RECT  0.9400 1.1750 1.0900 1.5700 ;
        RECT  0.7600 1.2800 1.0900 1.4000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5000 1.4650 3.7000 1.7250 ;
        RECT  0.5000 1.6900 3.6700 1.8100 ;
        RECT  3.5000 1.2200 3.6200 1.8100 ;
        RECT  0.5000 1.2200 0.6200 1.8100 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.0800 1.4100 6.2000 2.2100 ;
        RECT  4.4000 1.4100 6.2000 1.5300 ;
        RECT  5.6400 0.7950 5.9400 0.9150 ;
        RECT  5.8200 0.4000 5.9400 0.9150 ;
        RECT  4.0800 0.9300 5.7600 1.0500 ;
        RECT  5.6400 0.7950 5.7600 1.0500 ;
        RECT  5.2400 1.4100 5.3600 2.2100 ;
        RECT  5.0000 1.1750 5.1500 1.5300 ;
        RECT  5.0000 0.9300 5.1200 1.5300 ;
        RECT  4.9800 0.4000 5.1000 1.0500 ;
        RECT  4.4000 1.4100 4.5200 2.2100 ;
        RECT  4.0800 0.4000 4.2000 1.0500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.3800 0.1800 ;
        RECT  5.4000 -0.1800 5.5200 0.8100 ;
        RECT  4.5600 -0.1800 4.6800 0.8100 ;
        RECT  3.6000 0.4600 3.8400 0.5800 ;
        RECT  3.6000 -0.1800 3.7200 0.5800 ;
        RECT  0.3400 -0.1800 0.4600 0.6400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.3800 2.7900 ;
        RECT  5.6600 1.6500 5.7800 2.7900 ;
        RECT  4.8200 1.6500 4.9400 2.7900 ;
        RECT  3.8600 2.1700 4.1000 2.2900 ;
        RECT  3.8600 2.1700 3.9800 2.7900 ;
        RECT  2.9000 2.1700 3.1400 2.2900 ;
        RECT  2.9000 2.1700 3.0200 2.7900 ;
        RECT  1.9400 2.1700 2.1800 2.2900 ;
        RECT  1.9400 2.1700 2.0600 2.7900 ;
        RECT  0.9800 2.1700 1.2200 2.2900 ;
        RECT  0.9800 2.1700 1.1000 2.7900 ;
        RECT  0.1400 1.5600 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.8800 1.2900 3.9400 1.2900 3.9400 2.0500 3.5600 2.0500 3.5600 2.2100 3.4400 2.2100
                 3.4400 2.0500 2.6000 2.0500 2.6000 2.2100 2.4800 2.2100 2.4800 2.0500 1.6400 2.0500
                 1.6400 2.2100 1.5200 2.2100 1.5200 2.0500 0.6800 2.0500 0.6800 2.2100 0.5600 2.2100
                 0.5600 1.9300 3.8200 1.9300 3.8200 0.8200 2.2400 0.8200 2.2400 0.7700 2.1200 0.7700
                 2.1200 0.6500 2.3600 0.6500 2.3600 0.7000 3.9400 0.7000 3.9400 1.1700 4.8800 1.1700 ;
    END
END AND4X6

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.7700 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3500 0.7800 0.5300 1.1600 ;
        RECT  0.3300 0.7900 0.4800 1.1800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.7800 0.8200 1.2000 ;
        RECT  0.6500 0.7800 0.8200 1.1850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1350 0.9600 1.2550 1.2000 ;
        RECT  0.9400 0.9600 1.2550 1.1450 ;
        RECT  0.9400 0.8850 1.0900 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.4650 1.9600 1.7250 ;
        RECT  1.6750 1.3600 1.9300 1.4800 ;
        RECT  1.6750 1.2400 1.7950 1.4800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.0550 0.8850 3.4100 1.1450 ;
        RECT  3.0750 1.3200 3.1950 2.2100 ;
        RECT  3.0550 0.6800 3.1750 1.4400 ;
        RECT  2.2350 1.3200 3.1950 1.4400 ;
        RECT  2.0950 0.7300 3.1750 0.8500 ;
        RECT  2.8150 0.6800 3.1750 0.8500 ;
        RECT  2.2350 1.3200 2.3550 2.2100 ;
        RECT  1.9750 0.6800 2.2150 0.8000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.7700 0.1800 ;
        RECT  3.2950 -0.1800 3.4150 0.6700 ;
        RECT  2.3950 0.4900 2.6350 0.6100 ;
        RECT  2.3950 -0.1800 2.5150 0.6100 ;
        RECT  1.6150 -0.1800 1.7350 0.6700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.7700 2.7900 ;
        RECT  3.4950 1.5600 3.6150 2.7900 ;
        RECT  2.6550 1.5600 2.7750 2.7900 ;
        RECT  1.8150 1.8450 1.9350 2.7900 ;
        RECT  0.9750 1.5600 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.9350 1.1400 2.6950 1.1400 2.6950 1.1200 2.4750 1.1200 2.4750 1.1400 2.2350 1.1400
                 2.2350 1.1200 1.4950 1.1200 1.4950 1.3200 1.5150 1.3200 1.5150 2.2100 1.3950 2.2100
                 1.3950 1.4400 0.6750 1.4400 0.6750 2.2100 0.5550 2.2100 0.5550 1.3200 1.3750 1.3200
                 1.3750 0.6600 0.1600 0.6600 0.1600 0.5400 1.4950 0.5400 1.4950 1.0000 2.8150 1.0000
                 2.8150 1.0200 2.9350 1.0200 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.9000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3050 1.2250 0.5650 1.4950 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1750 1.0900 1.4400 ;
        RECT  0.8050 1.1750 1.0900 1.3450 ;
        RECT  0.8050 1.1000 0.9250 1.3450 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2250 1.0150 1.3800 1.4700 ;
        RECT  1.2250 1.0150 1.3450 1.4950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1050 1.9600 1.4350 ;
        RECT  1.7400 1.0900 1.8600 1.4150 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3200 0.8850 2.5400 1.1450 ;
        RECT  2.3200 0.6100 2.4400 1.4800 ;
        RECT  2.2250 1.3600 2.3450 2.0800 ;
        RECT  2.2200 0.4900 2.3400 0.7300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.9000 0.1800 ;
        RECT  2.6400 -0.1800 2.7600 0.7300 ;
        RECT  1.8000 -0.1800 1.9200 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.9000 2.7900 ;
        RECT  2.6450 1.4300 2.7650 2.7900 ;
        RECT  1.8050 1.5550 1.9250 2.7900 ;
        RECT  1.0250 2.1950 1.1450 2.7900 ;
        RECT  0.1350 2.1950 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2000 1.2400 2.0800 1.2400 2.0800 0.9700 1.6200 0.9700 1.6200 1.7350 1.5050 1.7350
                 1.5050 1.8550 1.3850 1.8550 1.3850 1.7350 0.4850 1.7350 0.4850 1.6150 1.5000 1.6150
                 1.5000 0.8600 0.2650 0.8600 0.2650 0.7400 1.6200 0.7400 1.6200 0.8500 2.2000 0.8500 ;
    END
END AND4X2

MACRO AND4X1
    CLASS CORE ;
    FOREIGN AND4X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0650 0.5100 1.4600 ;
        RECT  0.2400 1.0900 0.5100 1.2950 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7000 0.9300 0.8200 1.3550 ;
        RECT  0.6500 1.0550 0.8000 1.4600 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.0400 0.9300 1.1600 1.2800 ;
        RECT  0.9400 1.1100 1.0900 1.4600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5750 1.0200 1.6950 1.4600 ;
        RECT  1.5200 1.0200 1.6950 1.4400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3550 1.3400 2.4750 1.9900 ;
        RECT  2.0450 1.2300 2.4350 1.3800 ;
        RECT  2.3150 0.7300 2.4350 1.4600 ;
        RECT  2.2150 0.6100 2.3350 0.8500 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  1.7950 -0.1800 1.9150 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  1.9350 1.5000 2.0550 2.7900 ;
        RECT  1.0350 2.1400 1.1550 2.7900 ;
        RECT  0.1350 1.6200 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.1950 1.1100 1.9550 1.1100 1.9550 0.9000 1.4000 0.9000 1.4000 1.5800 1.6350 1.5800
                 1.6350 1.8200 1.5150 1.8200 1.5150 1.7000 0.4950 1.7000 0.4950 1.5800 1.2800 1.5800
                 1.2800 0.8100 0.2800 0.8100 0.2800 0.7900 0.1600 0.7900 0.1600 0.6700 0.4000 0.6700
                 0.4000 0.6900 1.4000 0.6900 1.4000 0.7800 2.0750 0.7800 2.0750 0.9900 2.1950 0.9900 ;
    END
END AND4X1

MACRO AND3XL
    CLASS CORE ;
    FOREIGN AND3XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3600 1.0400 0.5100 1.5000 ;
        RECT  0.3600 1.0400 0.4800 1.5300 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7700 1.0400 0.8900 1.3500 ;
        RECT  0.6500 1.1200 0.8000 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.2500 1.4650 1.6700 1.5850 ;
        RECT  1.2500 1.3450 1.3700 1.5850 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 1.1750 1.9600 1.4350 ;
        RECT  1.8300 1.1750 1.9500 2.0100 ;
        RECT  1.8100 0.6800 1.9300 1.4350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3900 -0.1800 1.5100 0.9200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.4100 1.8900 1.5300 2.7900 ;
        RECT  0.5700 1.8900 0.6900 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6900 1.3400 1.5700 1.3400 1.5700 1.2250 1.1300 1.2250 1.1300 1.8250 1.1100 1.8250
                 1.1100 2.0100 0.9900 2.0100 0.9900 1.7700 0.3300 1.7700 0.3300 1.9500 0.0900 1.9500
                 0.0900 1.8300 0.2100 1.8300 0.2100 1.6500 1.0100 1.6500 1.0100 0.9200 0.2900 0.9200
                 0.2900 0.6800 0.4100 0.6800 0.4100 0.8000 1.1300 0.8000 1.1300 1.1050 1.5700 1.1050
                 1.5700 1.1000 1.6900 1.1000 ;
    END
END AND3XL

MACRO AND3X8
    CLASS CORE ;
    FOREIGN AND3X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 6.0900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.4200 0.7500 2.5400 1.2200 ;
        RECT  0.3900 0.7500 2.5400 0.8700 ;
        RECT  0.4200 0.7500 0.5400 1.2200 ;
        RECT  0.3600 0.8850 0.5400 1.1450 ;
        RECT  0.3900 0.7500 0.5400 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.1750 2.2500 1.4350 ;
        RECT  2.1000 0.9900 2.2200 1.4350 ;
        RECT  1.2250 0.9900 2.2200 1.1100 ;
        RECT  0.9800 1.0400 1.3450 1.1600 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4650 1.2300 1.7250 1.5000 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.6400 0.7150 5.8800 0.8350 ;
        RECT  5.7200 1.2950 5.8400 2.2100 ;
        RECT  3.1800 0.7650 5.7600 0.8850 ;
        RECT  3.2000 1.2950 5.8400 1.4150 ;
        RECT  4.9000 0.7650 5.1500 1.1450 ;
        RECT  4.8000 0.7150 5.0400 0.8850 ;
        RECT  4.9000 0.7150 5.0200 1.4150 ;
        RECT  4.8800 1.2950 5.0000 2.2100 ;
        RECT  3.9600 0.7150 4.2000 0.8850 ;
        RECT  4.0400 1.2950 4.1600 2.2100 ;
        RECT  3.2000 1.2950 3.3200 2.2100 ;
        RECT  3.0600 0.7150 3.3000 0.8350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 6.0900 0.1800 ;
        RECT  5.2800 -0.1800 5.4000 0.6450 ;
        RECT  4.4400 -0.1800 4.5600 0.6450 ;
        RECT  3.5400 -0.1800 3.6600 0.6400 ;
        RECT  2.5800 -0.1800 2.8200 0.3900 ;
        RECT  0.5000 0.5100 0.7400 0.6300 ;
        RECT  0.5000 -0.1800 0.6200 0.6300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 6.0900 2.7900 ;
        RECT  5.3000 1.5350 5.4200 2.7900 ;
        RECT  4.4600 1.5350 4.5800 2.7900 ;
        RECT  3.6200 1.5350 3.7400 2.7900 ;
        RECT  2.7800 1.8600 2.9000 2.7900 ;
        RECT  1.9400 1.8600 2.0600 2.7900 ;
        RECT  1.1000 1.8600 1.2200 2.7900 ;
        RECT  0.2600 1.5600 0.3800 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.7800 1.1750 2.7800 1.1750 2.7800 1.7400 2.4800 1.7400 2.4800 2.2100 2.3600 2.2100
                 2.3600 1.7400 1.6400 1.7400 1.6400 2.2100 1.5200 2.2100 1.5200 1.7400 0.8000 1.7400
                 0.8000 2.2100 0.6800 2.2100 0.6800 1.5600 0.8000 1.5600 0.8000 1.6200 2.3600 1.6200
                 2.3600 1.5600 2.4800 1.5600 2.4800 1.6200 2.6600 1.6200 2.6600 0.6300 1.5600 0.6300
                 1.5600 0.5100 2.7800 0.5100 2.7800 1.0550 4.7800 1.0550 ;
    END
END AND3X8

MACRO AND3X6
    CLASS CORE ;
    FOREIGN AND3X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.2950 0.7500 2.4150 1.2200 ;
        RECT  0.3900 0.7500 2.4150 0.8700 ;
        RECT  0.4950 0.7500 0.6150 1.2200 ;
        RECT  0.3600 0.8850 0.6150 1.1450 ;
        RECT  0.3900 0.7500 0.6150 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.9900 2.0950 1.2300 ;
        RECT  1.8100 0.9900 1.9600 1.4350 ;
        RECT  0.9350 0.9900 2.0950 1.1100 ;
        RECT  0.7550 1.0400 1.0550 1.1600 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.2500 1.5550 1.5000 ;
        RECT  1.1750 1.2300 1.4350 1.5000 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.7550 1.3900 4.8750 2.2100 ;
        RECT  4.7350 0.4000 4.8550 0.9150 ;
        RECT  3.0750 1.3900 4.8750 1.5100 ;
        RECT  4.5550 0.7950 4.8550 0.9150 ;
        RECT  2.9950 0.9100 4.6750 1.0300 ;
        RECT  3.9550 1.1750 4.2800 1.5100 ;
        RECT  3.9550 0.9100 4.0750 1.5100 ;
        RECT  3.9150 1.3900 4.0350 2.2100 ;
        RECT  3.8950 0.4000 4.0150 1.0300 ;
        RECT  3.0750 1.3900 3.1950 2.2100 ;
        RECT  2.9950 0.4000 3.1150 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  4.3150 -0.1800 4.4350 0.7900 ;
        RECT  3.4750 -0.1800 3.5950 0.7900 ;
        RECT  2.4550 -0.1800 2.6950 0.3900 ;
        RECT  0.2750 0.5100 0.5150 0.6300 ;
        RECT  0.2750 -0.1800 0.3950 0.6300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  4.3350 1.6300 4.4550 2.7900 ;
        RECT  3.4950 1.6300 3.6150 2.7900 ;
        RECT  2.6550 1.8600 2.7750 2.7900 ;
        RECT  1.8150 1.8600 1.9350 2.7900 ;
        RECT  0.9750 1.8600 1.0950 2.7900 ;
        RECT  0.1350 1.5600 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.8350 1.2700 2.6550 1.2700 2.6550 1.7400 2.3550 1.7400 2.3550 2.2100 2.2350 2.2100
                 2.2350 1.7400 1.5150 1.7400 1.5150 2.2100 1.3950 2.2100 1.3950 1.7400 0.6750 1.7400
                 0.6750 2.2100 0.5550 2.2100 0.5550 1.5600 0.6750 1.5600 0.6750 1.6200 2.2350 1.6200
                 2.2350 1.5600 2.3550 1.5600 2.3550 1.6200 2.5350 1.6200 2.5350 0.6300 1.4350 0.6300
                 1.4350 0.5100 2.6550 0.5100 2.6550 1.1500 3.8350 1.1500 ;
    END
END AND3X6

MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.4800 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.7200 0.5100 1.2000 ;
        RECT  0.3600 0.7200 0.5100 1.1750 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8700 0.9600 0.9900 1.2000 ;
        RECT  0.6500 0.9600 0.9900 1.1450 ;
        RECT  0.6500 0.8850 0.8000 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.5200 1.4650 1.6700 1.7250 ;
        RECT  1.3500 1.3600 1.6400 1.4800 ;
        RECT  1.3500 1.2400 1.4700 1.4800 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.7900 0.8850 3.1200 1.1450 ;
        RECT  1.9100 1.3200 2.9100 1.4400 ;
        RECT  2.7900 0.6700 2.9100 1.4400 ;
        RECT  2.7500 1.3200 2.8700 2.2100 ;
        RECT  1.8300 0.7200 2.9100 0.8400 ;
        RECT  2.5500 0.6700 2.9100 0.8400 ;
        RECT  1.9100 1.3200 2.0300 2.2100 ;
        RECT  1.7100 0.6700 1.9500 0.7900 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.4800 0.1800 ;
        RECT  3.0300 -0.1800 3.1500 0.6600 ;
        RECT  2.1300 0.4800 2.3700 0.6000 ;
        RECT  2.1300 -0.1800 2.2500 0.6000 ;
        RECT  1.3500 -0.1800 1.4700 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.4800 2.7900 ;
        RECT  3.1700 1.5600 3.2900 2.7900 ;
        RECT  2.3300 1.5600 2.4500 2.7900 ;
        RECT  1.4900 1.8450 1.6100 2.7900 ;
        RECT  0.6500 1.5600 0.7700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.6700 1.1300 2.4300 1.1300 2.4300 1.1200 2.2100 1.1200 2.2100 1.1300 1.9700 1.1300
                 1.9700 1.1200 1.2300 1.1200 1.2300 1.4400 1.1900 1.4400 1.1900 2.2100 1.0700 2.2100
                 1.0700 1.4400 0.3500 1.4400 0.3500 2.2100 0.2300 2.2100 0.2300 1.3200 1.1100 1.3200
                 1.1100 0.6000 0.3300 0.6000 0.3300 0.4800 1.2300 0.4800 1.2300 1.0000 2.5500 1.0000
                 2.5500 1.0100 2.6700 1.0100 ;
    END
END AND3X4

MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.6100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 0.9850 0.2400 1.4350 ;
        RECT  0.1200 0.9600 0.2400 1.4350 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6750 0.9600 0.7950 1.3950 ;
        RECT  0.3600 1.0200 0.7950 1.1400 ;
        RECT  0.3600 1.0200 0.5100 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1550 1.2300 1.4350 1.4600 ;
        RECT  1.1550 1.2300 1.2750 1.6400 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8100 0.8850 1.9600 1.1450 ;
        RECT  1.8150 0.8850 1.9350 2.0350 ;
        RECT  1.6350 0.8850 1.9600 1.0250 ;
        RECT  1.6350 0.6100 1.7550 1.0250 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.6100 0.1800 ;
        RECT  2.0550 -0.1800 2.1750 0.6600 ;
        RECT  1.2150 -0.1800 1.3350 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.6100 2.7900 ;
        RECT  2.2350 1.3850 2.3550 2.7900 ;
        RECT  1.3950 1.6750 1.5150 2.7900 ;
        RECT  0.5550 1.7950 0.6750 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.5150 1.1100 1.0350 1.1100 1.0350 1.7600 1.0950 1.7600 1.0950 2.0000 0.9750 2.0000
                 0.9750 1.8800 0.9150 1.8800 0.9150 1.6750 0.3150 1.6750 0.3150 1.8550 0.0750 1.8550
                 0.0750 1.7350 0.1950 1.7350 0.1950 1.5550 0.9150 1.5550 0.9150 0.8400 0.1950 0.8400
                 0.1950 0.6000 0.3150 0.6000 0.3150 0.7200 1.0350 0.7200 1.0350 0.9900 1.5150 0.9900 ;
    END
END AND3X2

MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.3200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.0600 0.2400 1.5150 ;
        RECT  0.1200 1.0400 0.2400 1.5150 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7500 1.0400 0.8700 1.3500 ;
        RECT  0.3600 1.1200 0.8700 1.2400 ;
        RECT  0.3600 1.1200 0.5100 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.2300 1.1200 1.3800 1.5750 ;
        RECT  1.2300 1.0900 1.3500 1.5750 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.9300 1.1450 2.0500 2.0100 ;
        RECT  1.8100 0.8850 1.9600 1.2650 ;
        RECT  1.8100 0.6800 1.9300 1.2650 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.3200 0.1800 ;
        RECT  1.3900 -0.1800 1.5100 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.3200 2.7900 ;
        RECT  1.5100 1.5750 1.6300 2.7900 ;
        RECT  0.6150 2.2150 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.6900 1.2600 1.5700 1.2600 1.5700 0.9700 1.1100 0.9700 1.1100 1.6950 1.2100 1.6950
                 1.2100 1.9350 1.0900 1.9350 1.0900 1.8150 0.9900 1.8150 0.9900 1.7550 0.0750 1.7550
                 0.0750 1.6350 0.9900 1.6350 0.9900 0.9200 0.2700 0.9200 0.2700 0.6800 0.3900 0.6800
                 0.3900 0.8000 1.1100 0.8000 1.1100 0.8500 1.6900 0.8500 ;
    END
END AND3X1

MACRO AND2XL
    CLASS CORE ;
    FOREIGN AND2XL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.0700 1.1750 0.4150 1.2950 ;
        RECT  0.2950 1.0550 0.4150 1.2950 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.4650 1.0900 1.8200 ;
        RECT  0.8150 1.4650 1.0900 1.6100 ;
        RECT  0.8150 1.2500 0.9350 1.6100 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4850 1.4350 1.6050 1.8300 ;
        RECT  1.3500 1.4350 1.6050 1.5550 ;
        RECT  1.2300 1.1750 1.4700 1.4350 ;
        RECT  1.3500 0.5300 1.4700 1.5550 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.9300 -0.1800 1.0500 0.7700 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  1.0050 2.2300 1.1250 2.7900 ;
        RECT  0.1350 1.7100 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1100 1.1300 0.6750 1.1300 0.6750 1.8300 0.5550 1.8300 0.5550 0.9350 0.2900 0.9350
                 0.2900 0.5300 0.4100 0.5300 0.4100 0.8150 0.6750 0.8150 0.6750 1.0100 0.9900 1.0100
                 0.9900 0.8900 1.1100 0.8900 ;
    END
END AND2XL

MACRO AND2X8
    CLASS CORE ;
    FOREIGN AND2X8 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6500 0.9400 1.7700 1.2350 ;
        RECT  0.5950 0.9400 1.7700 1.0600 ;
        RECT  0.6300 0.9400 0.8700 1.1750 ;
        RECT  0.5950 0.9400 0.8700 1.0900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1750 1.1800 1.4350 1.4500 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.5300  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.9500 1.2950 5.0700 2.2100 ;
        RECT  4.8100 0.7150 5.0500 0.8350 ;
        RECT  2.4300 1.2950 5.0700 1.4150 ;
        RECT  2.3500 0.7650 4.9300 0.8850 ;
        RECT  4.1300 0.7650 4.2800 1.1450 ;
        RECT  4.1300 0.7150 4.2500 1.4150 ;
        RECT  4.1100 1.2950 4.2300 2.2100 ;
        RECT  3.9700 0.7150 4.2500 0.8850 ;
        RECT  3.2700 1.2950 3.3900 2.2100 ;
        RECT  3.1300 0.7150 3.3700 0.8850 ;
        RECT  2.4300 1.2950 2.5500 2.2100 ;
        RECT  2.2300 0.7150 2.4700 0.8350 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.2200 0.1800 ;
        RECT  4.4500 -0.1800 4.5700 0.6450 ;
        RECT  3.6100 -0.1800 3.7300 0.6450 ;
        RECT  2.7100 -0.1800 2.8300 0.6400 ;
        RECT  1.8100 0.4600 2.0500 0.5800 ;
        RECT  1.8100 -0.1800 1.9300 0.5800 ;
        RECT  0.5300 -0.1800 0.6500 0.7050 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.2200 2.7900 ;
        RECT  4.5300 1.5350 4.6500 2.7900 ;
        RECT  3.6900 1.5350 3.8100 2.7900 ;
        RECT  2.8500 1.5350 2.9700 2.7900 ;
        RECT  2.0100 1.8100 2.1300 2.7900 ;
        RECT  1.1700 1.8100 1.2900 2.7900 ;
        RECT  0.3300 1.5600 0.4500 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.0100 1.1750 2.0100 1.1750 2.0100 1.6900 1.7100 1.6900 1.7100 2.2100 1.5900 2.2100
                 1.5900 1.6900 0.8700 1.6900 0.8700 2.2100 0.7500 2.2100 0.7500 1.5600 0.8700 1.5600
                 0.8700 1.5700 1.5900 1.5700 1.5900 1.5600 1.7100 1.5600 1.7100 1.5700 1.8900 1.5700
                 1.8900 0.8200 1.1100 0.8200 1.1100 0.7000 2.0100 0.7000 2.0100 1.0550 4.0100 1.0550 ;
    END
END AND2X8

MACRO AND2X6
    CLASS CORE ;
    FOREIGN AND2X6 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.3500 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.6000 0.9400 1.7200 1.2600 ;
        RECT  0.3050 0.9400 1.7200 1.0600 ;
        RECT  0.4450 0.9400 0.5650 1.2600 ;
        RECT  0.3050 0.9400 0.5650 1.0900 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2160  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.8850 1.1800 1.1600 1.4250 ;
        RECT  0.8850 1.1800 1.1450 1.4450 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.2237  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0600 1.3900 4.1800 2.2100 ;
        RECT  3.9800 0.4000 4.1000 0.9150 ;
        RECT  2.3800 1.3900 4.1800 1.5100 ;
        RECT  3.8000 0.7950 4.1000 0.9150 ;
        RECT  2.2400 0.9100 3.9200 1.0300 ;
        RECT  3.2600 1.1750 3.4100 1.5100 ;
        RECT  3.2600 0.9100 3.3800 1.5100 ;
        RECT  3.2200 1.3900 3.3400 2.2100 ;
        RECT  3.1400 0.4000 3.2600 1.0300 ;
        RECT  2.3800 1.3900 2.5000 2.2100 ;
        RECT  2.2400 0.4000 2.3600 1.0300 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.3500 0.1800 ;
        RECT  3.5600 -0.1800 3.6800 0.7900 ;
        RECT  2.7200 -0.1800 2.8400 0.7900 ;
        RECT  1.7600 0.4600 2.0000 0.5800 ;
        RECT  1.7600 -0.1800 1.8800 0.5800 ;
        RECT  0.4800 -0.1800 0.6000 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.3500 2.7900 ;
        RECT  3.6400 1.6300 3.7600 2.7900 ;
        RECT  2.8000 1.6300 2.9200 2.7900 ;
        RECT  1.9600 1.8050 2.0800 2.7900 ;
        RECT  1.1200 1.8050 1.2400 2.7900 ;
        RECT  0.2800 1.5600 0.4000 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  3.1400 1.2700 1.9600 1.2700 1.9600 1.6850 1.6600 1.6850 1.6600 2.2100 1.5400 2.2100
                 1.5400 1.6850 0.8200 1.6850 0.8200 2.2100 0.7000 2.2100 0.7000 1.5650 1.5400 1.5650
                 1.5400 1.5600 1.6600 1.5600 1.6600 1.5650 1.8400 1.5650 1.8400 0.8200 1.0600 0.8200
                 1.0600 0.7000 1.9600 0.7000 1.9600 1.1500 3.1400 1.1500 ;
    END
END AND2X6

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 3.1900 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.3900 0.9700 0.5100 1.2100 ;
        RECT  0.0700 0.9700 0.5100 1.0900 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1080  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.3300 1.0900 1.7250 ;
        RECT  0.9500 1.2400 1.0700 1.7250 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3900 0.8850 2.5400 1.1450 ;
        RECT  1.5100 1.3200 2.5100 1.4400 ;
        RECT  2.3900 0.7600 2.5100 1.4400 ;
        RECT  2.3500 1.3200 2.4700 2.2100 ;
        RECT  1.5700 0.7600 2.5100 0.8800 ;
        RECT  2.3500 0.6400 2.4700 0.8800 ;
        RECT  1.4500 0.7100 1.6900 0.8300 ;
        RECT  1.5100 1.3200 1.6300 2.2100 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 3.1900 0.1800 ;
        RECT  2.7700 -0.1800 2.8900 0.7000 ;
        RECT  1.8700 0.5200 2.1100 0.6400 ;
        RECT  1.8700 -0.1800 1.9900 0.6400 ;
        RECT  1.0900 -0.1800 1.2100 0.7000 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 3.1900 2.7900 ;
        RECT  2.7700 1.5600 2.8900 2.7900 ;
        RECT  1.9300 1.5600 2.0500 2.7900 ;
        RECT  1.0900 1.8450 1.2100 2.7900 ;
        RECT  0.2500 1.5600 0.3700 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  2.2700 1.1700 2.0300 1.1700 2.0300 1.1200 1.8500 1.1200 1.8500 1.1700 1.6100 1.1700
                 1.6100 1.1200 0.7900 1.1200 0.7900 2.2100 0.6700 2.2100 0.6700 0.8300 0.3900 0.8300
                 0.3900 0.7100 0.7900 0.7100 0.7900 1.0000 2.1500 1.0000 2.1500 1.0500 2.2700 1.0500 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 2.0300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 1.0900 0.2900 1.4200 ;
        RECT  0.0700 1.1050 0.2200 1.4350 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.7150 1.0800 0.8350 1.4700 ;
        RECT  0.6500 1.0800 0.8350 1.4600 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3550 0.8850 1.6700 1.1450 ;
        RECT  1.3550 0.6700 1.4750 2.0700 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 2.0300 0.1800 ;
        RECT  1.7750 -0.1800 1.8950 0.7200 ;
        RECT  0.9350 -0.1800 1.0550 0.7200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 2.0300 2.7900 ;
        RECT  1.7750 1.4200 1.8950 2.7900 ;
        RECT  0.9350 1.5900 1.0550 2.7900 ;
        RECT  0.1350 2.2300 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.1950 1.2300 1.0750 1.2300 1.0750 0.9600 0.5300 0.9600 0.5300 1.5900 0.6350 1.5900
                 0.6350 1.8300 0.5150 1.8300 0.5150 1.7100 0.4100 1.7100 0.4100 0.9600 0.2350 0.9600
                 0.2350 0.6700 0.3550 0.6700 0.3550 0.8400 1.1950 0.8400 ;
    END
END AND2X2

MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 1.7400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 1.2850 0.2900 1.6100 ;
        RECT  0.0700 1.1750 0.2200 1.5050 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.0600  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6500 1.0500 0.8150 1.5050 ;
        RECT  0.6950 1.0200 0.8150 1.5050 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.3950 1.3400 1.5150 1.9900 ;
        RECT  1.3550 0.6800 1.4750 1.4600 ;
        RECT  1.1750 0.6500 1.4350 0.8000 ;
        RECT  1.3150 0.5600 1.4350 0.8000 ;
        END
    END Y
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 1.7400 0.1800 ;
        RECT  0.8950 -0.1800 1.0150 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 1.7400 2.7900 ;
        RECT  0.9750 1.6250 1.0950 2.7900 ;
        RECT  0.1350 1.7450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  1.2350 1.1100 0.9350 1.1100 0.9350 0.9000 0.5300 0.9000 0.5300 1.6250 0.6750 1.6250
                 0.6750 1.8650 0.5550 1.8650 0.5550 1.7450 0.4100 1.7450 0.4100 0.9000 0.1950 0.9000
                 0.1950 0.6100 0.3150 0.6100 0.3150 0.7800 1.0550 0.7800 1.0550 0.9900 1.2350 0.9900 ;
    END
END AND2X1

MACRO ADDHXL
    CLASS CORE ;
    FOREIGN ADDHXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.3050 0.4000 2.5450 0.5200 ;
        RECT  1.8250 1.0200 2.4250 1.1400 ;
        RECT  2.3050 0.4000 2.4250 1.1400 ;
        RECT  1.8250 0.4050 1.9450 1.1400 ;
        RECT  0.8550 0.4050 1.9450 0.5250 ;
        RECT  0.6500 0.8850 0.9750 1.0450 ;
        RECT  0.8550 0.4050 0.9750 1.0450 ;
        RECT  0.7000 0.8850 0.8200 1.1650 ;
        RECT  0.6500 0.8850 0.8200 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.9400 1.1700 1.2250 1.4000 ;
        RECT  1.1050 1.1550 1.2250 1.4000 ;
        RECT  0.9400 1.1700 1.0900 1.4350 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1350 0.5850 0.2550 1.8300 ;
        RECT  0.0700 1.1750 0.2550 1.4350 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.4050 0.7800 4.5250 1.7000 ;
        RECT  4.3850 1.4650 4.5050 1.8200 ;
        RECT  4.3850 0.6600 4.5050 0.9000 ;
        RECT  4.1300 1.4650 4.5050 1.7250 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  3.9450 -0.1800 4.0650 0.3800 ;
        RECT  2.0650 -0.1800 2.1850 0.9000 ;
        RECT  0.4950 0.6450 0.7350 0.7650 ;
        RECT  0.6150 -0.1800 0.7350 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  3.9450 2.2200 4.0650 2.7900 ;
        RECT  2.1050 1.7600 2.3450 1.8800 ;
        RECT  2.1050 1.7600 2.2250 2.7900 ;
        RECT  1.4550 2.0900 1.5750 2.7900 ;
        RECT  0.6150 2.2300 0.7350 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.2850 1.1800 3.8250 1.1800 3.8250 1.6600 3.4250 1.6600 3.4250 1.7600 3.1850 1.7600
                 3.1850 1.6400 3.3050 1.6400 3.3050 1.5400 3.7050 1.5400 3.7050 1.1800 3.1850 1.1800
                 3.1850 0.9000 3.0050 0.9000 3.0050 0.6600 3.1250 0.6600 3.1250 0.7800 3.3050 0.7800
                 3.3050 1.0600 4.2850 1.0600 ;
        POLYGON  3.7850 0.5200 2.7850 0.5200 2.7850 0.7800 2.7050 0.7800 2.7050 0.9000 2.6650 0.9000
                 2.6650 1.2800 2.8250 1.2800 2.8250 1.8200 2.7050 1.8200 2.7050 1.4000 2.5450 1.4000
                 2.5450 0.7800 2.5850 0.7800 2.5850 0.6600 2.6650 0.6600 2.6650 0.4000 3.7850 0.4000 ;
        POLYGON  3.5850 1.4200 3.0650 1.4200 3.0650 2.0600 2.4650 2.0600 2.4650 1.6400 1.8650 1.6400
                 1.8650 1.8200 1.7450 1.8200 1.7450 1.3800 1.5850 1.3800 1.5850 0.6600 1.7050 0.6600
                 1.7050 1.2600 1.8650 1.2600 1.8650 1.5200 2.5850 1.5200 2.5850 1.9400 2.9450 1.9400
                 2.9450 1.1600 2.7850 1.1600 2.7850 1.0400 3.0650 1.0400 3.0650 1.3000 3.5850 1.3000 ;
        POLYGON  1.4650 1.6750 1.1550 1.6750 1.1550 1.7700 0.9150 1.7700 0.9150 1.6750 0.4150 1.6750
                 0.4150 1.2700 0.5350 1.2700 0.5350 1.5550 1.3450 1.5550 1.3450 0.7650 1.1350 0.7650
                 1.1350 0.6450 1.4650 0.6450 ;
    END
END ADDHXL

MACRO ADDHX4
    CLASS CORE ;
    FOREIGN ADDHX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.8300 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.9150 0.8100 3.1550 0.9300 ;
        RECT  2.9150 0.3600 3.0350 0.9300 ;
        RECT  2.0750 0.3600 3.0350 0.4800 ;
        RECT  1.5950 0.9000 2.1950 1.0200 ;
        RECT  2.0750 0.3600 2.1950 1.0200 ;
        RECT  1.5950 0.3700 1.7150 1.0200 ;
        RECT  1.1150 0.3700 1.7150 0.4900 ;
        RECT  1.1150 0.3700 1.2350 0.9000 ;
        RECT  0.7550 0.7800 1.2350 0.9000 ;
        RECT  0.7550 0.7800 0.8750 1.1700 ;
        RECT  0.6500 0.8850 0.8750 1.1450 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2760  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.7350 1.7000 7.1350 1.8200 ;
        RECT  7.0150 1.0200 7.1350 1.8200 ;
        RECT  4.6750 1.9700 5.8550 2.0900 ;
        RECT  5.7350 1.7000 5.8550 2.0900 ;
        RECT  3.3500 2.1300 4.7950 2.2500 ;
        RECT  4.6750 1.9700 4.7950 2.2500 ;
        RECT  3.2750 1.0100 3.5150 1.1300 ;
        RECT  3.3500 1.0100 3.4700 2.2500 ;
        RECT  2.8350 1.3300 3.4700 1.4500 ;
        RECT  1.5100 1.7900 2.9550 1.9100 ;
        RECT  2.8350 1.3300 2.9550 1.9100 ;
        RECT  0.1700 1.7000 1.6300 1.8200 ;
        RECT  0.1700 1.0200 0.2900 1.8200 ;
        RECT  0.0700 1.1750 0.2900 1.4350 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.1000 1.5500 2.7150 1.6700 ;
        RECT  1.3550 1.1400 2.4350 1.2600 ;
        RECT  2.3150 0.6000 2.4350 1.2600 ;
        RECT  2.1000 1.1400 2.2500 1.6700 ;
        RECT  1.5150 1.4000 2.2500 1.5200 ;
        RECT  1.5150 1.4000 1.7550 1.5800 ;
        RECT  1.3550 0.6100 1.4750 1.2600 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4550 1.2200 6.5750 1.5800 ;
        RECT  5.3750 0.7400 6.5750 0.8600 ;
        RECT  5.4950 1.2200 6.5750 1.3400 ;
        RECT  6.1600 1.1750 6.3100 1.4350 ;
        RECT  6.1900 0.7400 6.3100 1.4350 ;
        RECT  5.4950 1.2200 5.6150 1.8500 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.8300 0.1800 ;
        RECT  6.8150 -0.1800 7.0550 0.3800 ;
        RECT  5.9150 -0.1800 6.0350 0.3800 ;
        RECT  4.8950 -0.1800 5.1350 0.3800 ;
        RECT  3.1550 -0.1800 3.2750 0.6500 ;
        RECT  1.8350 -0.1800 1.9550 0.7800 ;
        RECT  0.8750 -0.1800 0.9950 0.6600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.8300 2.7900 ;
        RECT  6.9350 1.9800 7.0550 2.7900 ;
        RECT  5.9750 1.9400 6.0950 2.7900 ;
        RECT  5.0150 2.2100 5.1350 2.7900 ;
        RECT  3.0750 1.5700 3.1950 2.7900 ;
        RECT  1.9950 2.0300 2.2350 2.7900 ;
        RECT  1.0350 1.9400 1.2750 2.7900 ;
        RECT  0.1350 1.9400 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.4750 1.4600 7.4150 1.4600 7.4150 1.5800 7.2950 1.5800 7.2950 1.3400 7.3550 1.3400
                 7.3550 0.6200 4.6550 0.6200 4.6550 0.5300 4.0750 0.5300 4.0750 0.9100 4.2550 0.9100
                 4.2550 1.1100 4.5750 1.1100 4.5750 1.3700 4.4550 1.3700 4.4550 1.2300 4.1350 1.2300
                 4.1350 1.1500 3.8750 1.1500 3.8750 0.9100 3.9550 0.9100 3.9550 0.4100 4.7750 0.4100
                 4.7750 0.5000 7.3550 0.5000 7.3550 0.4900 7.4750 0.4900 ;
        POLYGON  5.2550 1.2400 5.1550 1.2400 5.1550 1.8500 4.4950 1.8500 4.4950 2.0100 4.2550 2.0100
                 4.2550 1.7300 5.0350 1.7300 5.0350 0.9900 4.3750 0.9900 4.3750 0.7700 4.1950 0.7700
                 4.1950 0.6500 4.4950 0.6500 4.4950 0.8700 5.2550 0.8700 ;
        POLYGON  4.9150 1.6100 4.0150 1.6100 4.0150 1.8500 3.8950 1.8500 3.8950 1.3900 3.6350 1.3900
                 3.6350 0.6700 3.7150 0.6700 3.7150 0.4100 3.8350 0.4100 3.8350 0.7900 3.7550 0.7900
                 3.7550 1.2700 4.0150 1.2700 4.0150 1.4900 4.7950 1.4900 4.7950 1.1100 4.9150 1.1100 ;
        POLYGON  1.2350 1.4100 0.7350 1.4100 0.7350 1.5800 0.6150 1.5800 0.6150 1.4100 0.4100 1.4100
                 0.4100 0.9000 0.2350 0.9000 0.2350 0.6100 0.3550 0.6100 0.3550 0.7800 0.5300 0.7800
                 0.5300 1.2900 1.1150 1.2900 1.1150 1.0200 1.2350 1.0200 ;
    END
END ADDHX4

MACRO ADDHX2
    CLASS CORE ;
    FOREIGN ADDHX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.5100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0750 0.4200 5.3150 0.5400 ;
        RECT  3.4850 0.5000 5.1950 0.6200 ;
        RECT  1.2550 0.4800 3.6050 0.6000 ;
        RECT  3.2150 0.3800 3.4550 0.6000 ;
        RECT  2.8150 0.4800 2.9350 1.4600 ;
        RECT  0.5350 0.6450 1.3750 0.7650 ;
        RECT  1.2550 0.4800 1.3750 0.7650 ;
        RECT  0.5350 0.8850 0.8000 1.1450 ;
        RECT  0.5350 0.6450 0.6550 1.2400 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5400 1.9400 2.6600 2.2400 ;
        RECT  2.3800 1.9400 2.6600 2.0600 ;
        RECT  1.3150 1.8600 2.5000 1.9800 ;
        RECT  1.3150 1.3000 1.4350 1.9800 ;
        RECT  1.1750 1.3000 1.4350 1.6700 ;
        RECT  1.1600 1.3000 1.4350 1.4200 ;
        END
    END A
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.8000 1.4650 1.9600 1.7250 ;
        RECT  1.6600 1.6200 1.9200 1.7400 ;
        RECT  1.8000 0.7200 1.9200 1.7400 ;
        RECT  1.4950 0.7200 1.9200 0.8400 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3550 0.8850 4.5700 1.1450 ;
        RECT  4.3200 1.4000 4.5600 1.5200 ;
        RECT  4.3550 0.7400 4.4750 1.5200 ;
        RECT  4.2350 0.7400 4.4750 0.8600 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 5.5100 0.1800 ;
        RECT  4.7150 -0.1800 4.9550 0.3800 ;
        RECT  3.7550 -0.1800 3.9950 0.3800 ;
        RECT  1.9750 -0.1800 2.2150 0.3600 ;
        RECT  1.0150 -0.1800 1.1350 0.3800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 5.5100 2.7900 ;
        RECT  4.8000 2.0400 5.0400 2.1600 ;
        RECT  4.8000 2.0400 4.9200 2.7900 ;
        RECT  3.8400 1.8800 4.0800 2.0000 ;
        RECT  3.8400 1.8800 3.9600 2.7900 ;
        RECT  2.2000 2.2200 2.3200 2.7900 ;
        RECT  1.1800 2.1000 1.4200 2.2200 ;
        RECT  1.1800 2.1000 1.3000 2.7900 ;
        RECT  0.3400 1.6800 0.4600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  5.4350 0.8600 5.3750 0.8600 5.3750 1.7600 3.9300 1.7600 3.9300 1.4800 3.2950 1.4800
                 3.2950 1.2400 3.4150 1.2400 3.4150 1.3600 4.0500 1.3600 4.0500 1.6400 5.2550 1.6400
                 5.2550 0.8600 5.1950 0.8600 5.1950 0.7400 5.4350 0.7400 ;
        POLYGON  4.2200 1.2400 4.1000 1.2400 4.1000 1.1200 3.1750 1.1200 3.1750 1.7000 3.1600 1.7000
                 3.1600 1.8200 3.0400 1.8200 3.0400 1.5800 3.0550 1.5800 3.0550 0.7200 3.2950 0.7200
                 3.2950 0.8400 3.1750 0.8400 3.1750 1.0000 4.2200 1.0000 ;
        POLYGON  3.7200 2.1800 2.7800 2.1800 2.7800 1.8200 2.6200 1.8200 2.6200 1.7000 2.5750 1.7000
                 2.5750 0.8400 2.4550 0.8400 2.4550 0.7200 2.6950 0.7200 2.6950 1.5800 2.7400 1.5800
                 2.7400 1.7000 2.9000 1.7000 2.9000 2.0600 3.7200 2.0600 ;
        POLYGON  1.6800 1.3000 1.5600 1.3000 1.5600 1.1800 1.0400 1.1800 1.0400 1.7400 0.7000 1.7400
                 0.7000 1.6200 0.9200 1.6200 0.9200 1.4800 0.2950 1.4800 0.2950 0.6600 0.4150 0.6600
                 0.4150 1.3600 0.9200 1.3600 0.9200 1.0600 1.6800 1.0600 ;
    END
END ADDHX2

MACRO ADDHX1
    CLASS CORE ;
    FOREIGN ADDHX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 4.6400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1200  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  2.5200 0.3600 2.8000 0.4800 ;
        RECT  2.0400 0.6500 2.6400 0.7700 ;
        RECT  2.5200 0.3600 2.6400 0.7700 ;
        RECT  2.0400 0.3800 2.1600 0.7700 ;
        RECT  0.8900 0.3800 2.1600 0.5000 ;
        RECT  0.7350 0.7100 1.0100 0.8300 ;
        RECT  0.8900 0.3800 1.0100 0.8300 ;
        RECT  0.7300 0.9800 0.9700 1.1000 ;
        RECT  0.5950 0.9400 0.8550 1.0900 ;
        RECT  0.7350 0.7100 0.8550 1.1000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.1400 0.9000 1.4350 1.1350 ;
        RECT  1.1300 0.9000 1.4350 1.1100 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1700 0.6000 0.2900 2.2100 ;
        RECT  0.0700 1.1750 0.2900 1.4350 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.3800 1.1750 4.5700 1.4350 ;
        RECT  4.3800 0.8000 4.5000 1.4350 ;
        RECT  4.3600 1.3000 4.4800 1.9900 ;
        RECT  4.3600 0.6800 4.4800 0.9200 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 4.6400 0.1800 ;
        RECT  3.8800 0.6800 4.1200 0.8000 ;
        RECT  3.9800 -0.1800 4.1000 0.8000 ;
        RECT  2.2800 -0.1800 2.4000 0.5300 ;
        RECT  0.5300 0.4700 0.7700 0.5900 ;
        RECT  0.6500 -0.1800 0.7700 0.5900 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 4.6400 2.7900 ;
        RECT  3.9400 1.7200 4.0600 2.7900 ;
        RECT  2.2200 1.8500 2.4600 1.9700 ;
        RECT  2.2200 1.8500 2.3400 2.7900 ;
        RECT  1.4900 2.0200 1.6100 2.7900 ;
        RECT  0.5300 1.9100 0.7700 2.1500 ;
        RECT  0.5300 1.9100 0.6500 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  4.2600 1.1800 4.0200 1.1800 4.0200 1.1200 3.8800 1.1200 3.8800 1.6000 3.4200 1.6000
                 3.4200 1.8700 3.3000 1.8700 3.3000 1.4800 3.7600 1.4800 3.7600 1.1200 3.3000 1.1200
                 3.3000 0.8600 3.1800 0.8600 3.1800 0.6200 3.3000 0.6200 3.3000 0.7400 3.4200 0.7400
                 3.4200 1.0000 4.1400 1.0000 4.1400 1.0600 4.2600 1.0600 ;
        POLYGON  3.8600 0.4800 3.7400 0.4800 3.7400 0.5000 3.0400 0.5000 3.0400 0.7400 2.8800 0.7400
                 2.8800 1.0100 2.7400 1.0100 2.7400 1.3700 2.9400 1.3700 2.9400 1.8700 2.8200 1.8700
                 2.8200 1.4900 2.6200 1.4900 2.6200 0.8900 2.7600 0.8900 2.7600 0.6200 2.9200 0.6200
                 2.9200 0.3800 3.6200 0.3800 3.6200 0.3600 3.8600 0.3600 ;
        POLYGON  3.6400 1.3600 3.1800 1.3600 3.1800 2.1100 2.5800 2.1100 2.5800 1.7300 1.9200 1.7300
                 1.9200 1.8700 1.8000 1.8700 1.8000 0.6200 1.9200 0.6200 1.9200 1.6100 2.7000 1.6100
                 2.7000 1.9900 3.0600 1.9900 3.0600 1.2500 2.8600 1.2500 2.8600 1.1300 3.1800 1.1300
                 3.1800 1.2400 3.6400 1.2400 ;
        POLYGON  1.6750 1.3750 1.1300 1.3750 1.1300 2.0900 1.0100 2.0900 1.0100 1.3750 0.5700 1.3750
                 0.5700 1.4800 0.4500 1.4800 0.4500 1.2400 0.5700 1.2400 0.5700 1.2550 1.5550 1.2550
                 1.5550 0.7800 1.2300 0.7800 1.2300 0.6600 1.6750 0.6600 ;
    END
END ADDHX1

MACRO ADDFXL
    CLASS CORE ;
    FOREIGN ADDFXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.2350 0.7800 5.9700 0.9000 ;
        RECT  2.6250 0.7200 3.3550 0.8000 ;
        RECT  2.7050 0.7800 5.9700 0.8400 ;
        RECT  2.6250 0.6500 2.8850 0.8000 ;
        RECT  2.7050 0.6500 2.8250 0.9600 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4900 1.0200 6.6100 1.5000 ;
        RECT  6.4500 1.0200 6.6100 1.4350 ;
        RECT  2.0450 1.0800 6.6100 1.1400 ;
        RECT  3.5850 1.0200 6.6100 1.1400 ;
        RECT  2.2600 1.0800 3.7050 1.2000 ;
        RECT  1.4450 1.0200 2.3800 1.0800 ;
        RECT  1.4450 0.9600 2.1650 1.0800 ;
        RECT  1.3250 1.0800 1.5650 1.2000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.9750 1.2600 6.3300 1.3800 ;
        RECT  1.8050 1.3200 4.0950 1.4400 ;
        RECT  2.9150 1.3200 3.1750 1.6700 ;
        RECT  1.8050 1.2000 1.9250 1.4400 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5550 1.6050 0.6750 1.9650 ;
        RECT  0.1550 1.0050 0.6750 1.1250 ;
        RECT  0.5550 0.6450 0.6750 1.1250 ;
        RECT  0.0700 1.6050 0.6750 1.7250 ;
        RECT  0.0700 1.4650 0.2750 1.7250 ;
        RECT  0.1550 1.0050 0.2750 1.7250 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.1680  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.1750 0.4000 7.2950 0.6400 ;
        RECT  7.0300 1.4650 7.1800 1.7250 ;
        RECT  7.0550 0.5200 7.1750 1.7250 ;
        RECT  7.0500 1.4650 7.1700 2.0900 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.7550 -0.1800 6.8750 0.6400 ;
        RECT  4.5450 0.3000 4.7850 0.4200 ;
        RECT  4.5450 -0.1800 4.6650 0.4200 ;
        RECT  3.7050 -0.1800 3.8250 0.6400 ;
        RECT  1.5450 -0.1800 1.7850 0.3200 ;
        RECT  0.1350 -0.1800 0.2550 0.8850 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.5700 1.9800 6.6900 2.7900 ;
        RECT  4.0600 2.2200 4.3000 2.7900 ;
        RECT  3.5200 2.1600 3.6400 2.7900 ;
        RECT  1.4250 2.0400 1.5450 2.7900 ;
        RECT  0.1350 1.8450 0.2550 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  6.9350 1.3450 6.8500 1.3450 6.8500 1.8600 5.8300 1.8600 5.8300 2.0300 5.5900 2.0300
                 5.5900 1.8600 5.3800 1.8600 5.3800 2.0000 5.2600 2.0000 5.2600 1.7400 6.7300 1.7400
                 6.7300 0.8800 6.5150 0.8800 6.5150 0.5800 5.4450 0.5800 5.4450 0.4600 6.6350 0.4600
                 6.6350 0.7600 6.8500 0.7600 6.8500 1.1050 6.9350 1.1050 ;
        POLYGON  5.2650 0.5800 5.1450 0.5800 5.1450 0.6600 4.1850 0.6600 4.1850 0.5800 4.0650 0.5800
                 4.0650 0.4600 4.3050 0.4600 4.3050 0.5400 5.0250 0.5400 5.0250 0.4600 5.2650 0.4600 ;
        POLYGON  5.1600 1.6200 5.1400 1.6200 5.1400 2.1800 4.4200 2.1800 4.4200 2.1000 3.8500 2.1000
                 3.8500 2.0400 3.5850 2.0400 3.5850 2.0300 2.7900 2.0300 2.7900 1.9600 1.6650 1.9600
                 1.6650 1.9200 0.8250 1.9200 0.8250 1.3650 0.5150 1.3650 0.5150 1.4850 0.3950 1.4850
                 0.3950 1.2450 0.8250 1.2450 0.8250 0.4400 2.3850 0.4400 2.3850 0.4100 3.1250 0.4100
                 3.1250 0.4600 3.2450 0.4600 3.2450 0.5800 3.0050 0.5800 3.0050 0.5300 2.5050 0.5300
                 2.5050 0.9000 2.3850 0.9000 2.3850 0.5600 0.9450 0.5600 0.9450 1.8000 1.7850 1.8000
                 1.7850 1.8400 2.3850 1.8400 2.3850 1.6600 2.5050 1.6600 2.5050 1.8400 2.7900 1.8400
                 2.7900 1.7900 2.9100 1.7900 2.9100 1.9100 3.7050 1.9100 3.7050 1.9200 3.9700 1.9200
                 3.9700 1.9800 4.5400 1.9800 4.5400 2.0600 5.0200 2.0600 5.0200 1.6200 4.9200 1.6200
                 4.9200 1.5000 5.1600 1.5000 ;
        POLYGON  4.9000 1.9400 4.6600 1.9400 4.6600 1.8000 3.8800 1.8000 3.8800 1.5600 4.0000 1.5600
                 4.0000 1.6800 4.7800 1.6800 4.7800 1.8200 4.9000 1.8200 ;
        POLYGON  2.1450 0.8400 1.2450 0.8400 1.2450 0.9200 1.1250 0.9200 1.1250 0.6800 1.2450 0.6800
                 1.2450 0.7200 2.1450 0.7200 ;
        POLYGON  2.1450 1.7200 1.9050 1.7200 1.9050 1.6800 1.0650 1.6800 1.0650 1.5600 2.0250 1.5600
                 2.0250 1.6000 2.1450 1.6000 ;
    END
END ADDFXL

MACRO ADDFX4
    CLASS CORE ;
    FOREIGN ADDFX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3240  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0350 0.8200 7.4950 0.9400 ;
        RECT  5.1750 0.8200 5.4150 1.0900 ;
        RECT  4.0550 0.7800 5.1550 0.9000 ;
        RECT  4.0750 0.6500 4.3350 0.9000 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2750 0.9400 8.3950 1.2500 ;
        RECT  8.1350 0.9400 8.3950 1.1600 ;
        RECT  7.6550 1.0400 8.3950 1.1600 ;
        RECT  5.5350 1.0600 7.7750 1.1800 ;
        RECT  4.7950 1.2100 5.6550 1.3300 ;
        RECT  5.5350 1.0600 5.6550 1.3300 ;
        RECT  4.7950 1.0200 4.9150 1.3300 ;
        RECT  3.7350 1.0200 4.9150 1.1400 ;
        RECT  2.6750 0.9800 3.8550 1.1000 ;
        RECT  2.6750 0.9800 2.7950 1.2400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8950 1.2800 8.1350 1.4000 ;
        RECT  5.7750 1.3000 8.0150 1.4200 ;
        RECT  4.4200 1.4500 5.8950 1.5700 ;
        RECT  5.7750 1.3000 5.8950 1.5700 ;
        RECT  4.4200 1.2800 4.6750 1.5700 ;
        RECT  4.4200 1.2800 4.5700 1.7250 ;
        RECT  4.0500 1.2800 4.6750 1.4000 ;
        RECT  3.1350 1.2600 4.1700 1.3400 ;
        RECT  3.2550 1.2800 4.6750 1.3800 ;
        RECT  3.1350 1.2200 3.3750 1.3400 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4350 1.3200 1.5550 2.2100 ;
        RECT  1.4350 0.6700 1.5550 0.9600 ;
        RECT  0.5550 1.3200 1.5550 1.4400 ;
        RECT  0.5550 0.8400 1.5550 0.9600 ;
        RECT  0.5950 1.3200 0.7150 2.2100 ;
        RECT  0.5950 0.6700 0.7150 0.9600 ;
        RECT  0.5550 0.7900 0.6750 1.4400 ;
        RECT  0.3600 0.8850 0.6750 1.1450 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.7350 0.8850 10.0800 1.1450 ;
        RECT  8.8550 1.3200 9.8550 1.4400 ;
        RECT  9.7350 0.7600 9.8550 1.4400 ;
        RECT  9.6950 1.3200 9.8150 2.2100 ;
        RECT  8.8550 0.7600 9.8550 0.8800 ;
        RECT  9.6950 0.5900 9.8150 0.8800 ;
        RECT  8.8550 1.3200 8.9750 2.2100 ;
        RECT  8.8550 0.5900 8.9750 0.8800 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  10.1150 -0.1800 10.2350 0.6400 ;
        RECT  9.2750 -0.1800 9.3950 0.6400 ;
        RECT  8.3750 0.4600 8.6150 0.5800 ;
        RECT  8.3750 -0.1800 8.4950 0.5800 ;
        RECT  5.9350 0.3400 6.1750 0.4600 ;
        RECT  5.9350 -0.1800 6.0550 0.4600 ;
        RECT  5.0950 -0.1800 5.2150 0.6400 ;
        RECT  2.8150 -0.1800 3.0550 0.3800 ;
        RECT  1.8550 -0.1800 1.9750 0.7200 ;
        RECT  1.0150 -0.1800 1.1350 0.7200 ;
        RECT  0.1750 -0.1800 0.2950 0.7200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  10.1150 1.5600 10.2350 2.7900 ;
        RECT  9.2750 1.5600 9.3950 2.7900 ;
        RECT  8.3750 2.0200 8.6150 2.1500 ;
        RECT  8.3750 2.0200 8.4950 2.7900 ;
        RECT  5.9350 2.1700 6.1750 2.7900 ;
        RECT  4.9750 2.1700 5.2150 2.7900 ;
        RECT  2.8750 2.1000 2.9950 2.7900 ;
        RECT  1.7950 2.0300 2.0350 2.1500 ;
        RECT  1.7950 2.0300 1.9150 2.7900 ;
        RECT  1.0150 1.5600 1.1350 2.7900 ;
        RECT  0.1750 1.5600 0.2950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.6150 1.1200 8.6350 1.1200 8.6350 1.9000 7.6550 1.9000 7.6550 2.1500 7.4150 2.1500
                 7.4150 1.9000 7.2550 1.9000 7.2550 2.1500 7.0150 2.1500 7.0150 1.8800 7.1350 1.8800
                 7.1350 1.7800 8.5150 1.7800 8.5150 0.8200 8.1350 0.8200 8.1350 0.7000 6.8350 0.7000
                 6.8350 0.5800 7.5150 0.5800 7.5150 0.5000 7.7550 0.5000 7.7550 0.5800 8.2550 0.5800
                 8.2550 0.7000 8.6350 0.7000 8.6350 1.0000 9.6150 1.0000 ;
        POLYGON  7.3350 1.6600 6.8950 1.6600 6.8950 2.0500 4.4550 2.0500 4.4550 2.2100 4.3350 2.2100
                 4.3350 2.0500 3.8950 2.0500 3.8950 2.1500 3.7750 2.1500 3.7750 2.0500 3.6850 2.0500
                 3.6850 1.9800 2.3600 1.9800 2.3600 1.9100 2.0950 1.9100 2.0950 1.2000 0.7950 1.2000
                 0.7950 1.0800 2.0950 1.0800 2.0950 0.5000 3.7750 0.5000 3.7750 0.4100 4.5750 0.4100
                 4.5750 0.6500 4.4550 0.6500 4.4550 0.5300 3.8950 0.5300 3.8950 0.7400 3.7750 0.7400
                 3.7750 0.6200 2.2150 0.6200 2.2150 1.7900 2.4800 1.7900 2.4800 1.8600 3.7750 1.8600
                 3.7750 1.5000 3.8950 1.5000 3.8950 1.9300 4.3350 1.9300 4.3350 1.8450 4.4550 1.8450
                 4.4550 1.9300 6.7750 1.9300 6.7750 1.5400 7.3350 1.5400 ;
        RECT  5.4550 0.5800 6.6550 0.7000 ;
        POLYGON  6.6550 1.8100 5.4550 1.8100 5.4550 1.6900 6.4150 1.6900 6.4150 1.6200 6.6550 1.6200 ;
        RECT  2.3350 0.7400 3.5350 0.8600 ;
        POLYGON  3.4750 1.7400 3.3550 1.7400 3.3550 1.6200 2.5150 1.6200 2.5150 1.6700 2.3950 1.6700
                 2.3950 1.3400 2.5150 1.3400 2.5150 1.5000 3.4750 1.5000 ;
    END
END ADDFX4

MACRO ADDFX2
    CLASS CORE ;
    FOREIGN ADDFX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.4100 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0000 0.8300 6.5150 0.9500 ;
        RECT  3.1250 0.7600 4.1200 0.8800 ;
        RECT  3.2050 0.6500 3.4650 0.8800 ;
        RECT  3.1250 0.7100 3.2450 0.9500 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9750 1.0700 7.2350 1.3800 ;
        RECT  2.8750 1.0700 7.2350 1.1900 ;
        RECT  3.8150 1.0700 4.0550 1.2000 ;
        RECT  1.8650 1.0200 2.9950 1.1400 ;
        RECT  1.7450 1.0800 1.9850 1.2000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.6400 1.3100 6.8550 1.4300 ;
        RECT  2.6350 1.3200 4.8800 1.4400 ;
        RECT  3.5500 1.3200 3.7000 1.7250 ;
        RECT  3.2750 1.3100 3.5550 1.4400 ;
        RECT  2.1650 1.2600 2.7550 1.3800 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.6450 0.6800 0.7650 2.2100 ;
        RECT  0.3600 1.1750 0.7650 1.2950 ;
        RECT  0.3600 1.1750 0.5100 1.4350 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.6950 0.8850 8.0500 1.1450 ;
        RECT  7.6350 1.6200 7.8750 2.1500 ;
        RECT  7.6950 0.6400 7.8150 2.1500 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.4100 0.1800 ;
        RECT  8.1150 -0.1800 8.2350 0.6900 ;
        RECT  7.2750 -0.1800 7.3950 0.6900 ;
        RECT  5.0650 0.3500 5.3050 0.4700 ;
        RECT  5.0650 -0.1800 5.1850 0.4700 ;
        RECT  4.1650 0.4600 4.4050 0.5800 ;
        RECT  4.1650 -0.1800 4.2850 0.5800 ;
        RECT  1.9650 -0.1800 2.2050 0.3200 ;
        RECT  1.0650 -0.1800 1.1850 0.7300 ;
        RECT  0.2250 -0.1800 0.3450 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.4100 2.7900 ;
        RECT  8.1150 1.5600 8.2350 2.7900 ;
        RECT  7.2150 2.0300 7.4550 2.1500 ;
        RECT  7.2150 2.0300 7.3350 2.7900 ;
        RECT  4.6750 2.2700 4.9150 2.7900 ;
        RECT  3.8950 2.0850 4.0150 2.7900 ;
        RECT  1.8450 2.0000 1.9650 2.7900 ;
        RECT  1.0050 1.9800 1.2450 2.1500 ;
        RECT  1.0050 1.9800 1.1250 2.7900 ;
        RECT  0.2250 1.5600 0.3450 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.5550 1.3000 7.4750 1.3000 7.4750 1.9100 6.5350 1.9100 6.5350 2.0900 6.4150 2.0900
                 6.4150 1.9100 5.7550 1.9100 5.7550 1.7900 7.3550 1.7900 7.3550 0.9300 7.0350 0.9300
                 7.0350 0.6300 6.1450 0.6300 6.1450 0.6400 6.0250 0.6400 6.0250 0.4000 6.1450 0.4000
                 6.1450 0.5100 7.1550 0.5100 7.1550 0.8100 7.4750 0.8100 7.4750 1.0600 7.5550 1.0600 ;
        POLYGON  6.3150 1.6700 5.6350 1.6700 5.6350 2.0300 4.8400 2.0300 4.8400 2.0500 4.1350 2.0500
                 4.1350 1.9650 3.1950 1.9650 3.1950 1.9600 2.0850 1.9600 2.0850 1.8600 1.3050 1.8600
                 1.3050 1.2600 0.8850 1.2600 0.8850 1.1400 1.3050 1.1400 1.3050 0.4400 2.9650 0.4400
                 2.9650 0.4100 3.5850 0.4100 3.5850 0.4000 3.7050 0.4000 3.7050 0.6400 3.5850 0.6400
                 3.5850 0.5300 3.0850 0.5300 3.0850 0.5600 2.9250 0.5600 2.9250 0.9000 2.8050 0.9000
                 2.8050 0.5600 1.4250 0.5600 1.4250 1.7400 2.2050 1.7400 2.2050 1.8400 2.8050 1.8400
                 2.8050 1.6600 2.9250 1.6600 2.9250 1.8400 3.1950 1.8400 3.1950 1.6900 3.3150 1.6900
                 3.3150 1.8450 4.2550 1.8450 4.2550 1.9300 4.7200 1.9300 4.7200 1.9100 5.5150 1.9100
                 5.5150 1.5500 6.3150 1.5500 ;
        POLYGON  5.7850 0.5800 5.6650 0.5800 5.6650 0.7100 4.7050 0.7100 4.7050 0.5800 4.5850 0.5800
                 4.5850 0.4600 4.8250 0.4600 4.8250 0.5900 5.5450 0.5900 5.5450 0.4600 5.7850 0.4600 ;
        POLYGON  5.3950 1.7900 4.4950 1.7900 4.4950 1.8100 4.3750 1.8100 4.3750 1.5700 4.4950 1.5700
                 4.4950 1.6700 5.3950 1.6700 ;
        POLYGON  2.5650 0.8400 1.6650 0.8400 1.6650 0.9200 1.5450 0.9200 1.5450 0.6800 1.6650 0.6800
                 1.6650 0.7200 2.5650 0.7200 ;
        POLYGON  2.5650 1.7200 2.3250 1.7200 2.3250 1.6200 1.5450 1.6200 1.5450 1.3800 1.6650 1.3800
                 1.6650 1.5000 2.4450 1.5000 2.4450 1.6000 2.5650 1.6000 ;
    END
END ADDFX2

MACRO ADDFX1
    CLASS CORE ;
    FOREIGN ADDFX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 7.5400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1800  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.7650 0.8300 5.9900 0.9500 ;
        RECT  2.7050 0.7800 3.9650 0.8800 ;
        RECT  3.5000 0.8300 5.9900 0.9000 ;
        RECT  2.6250 0.7600 3.6200 0.8000 ;
        RECT  2.6250 0.6500 2.8850 0.8000 ;
        RECT  2.7050 0.6500 2.8250 0.9800 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.4500 1.0700 6.7350 1.2900 ;
        RECT  6.6150 1.0500 6.7350 1.2900 ;
        RECT  6.4500 1.0700 6.6000 1.4350 ;
        RECT  3.5500 1.0700 6.7350 1.1900 ;
        RECT  2.0650 1.1000 3.6700 1.2200 ;
        RECT  1.4650 0.9800 2.1850 1.1000 ;
        RECT  1.3450 1.0600 1.5850 1.1800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2400  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.8650 1.3100 6.3300 1.4300 ;
        RECT  1.8250 1.3400 3.9850 1.4600 ;
        RECT  3.2050 1.3400 3.4650 1.6700 ;
        RECT  1.8250 1.2200 1.9450 1.4600 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5600 1.3150 0.6800 2.2050 ;
        RECT  0.1000 0.8350 0.6800 0.9550 ;
        RECT  0.5600 0.6650 0.6800 0.9550 ;
        RECT  0.0700 1.3150 0.6800 1.4350 ;
        RECT  0.0700 1.1750 0.2200 1.4350 ;
        RECT  0.1000 0.8350 0.2200 1.4350 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.2750 0.8850 7.4700 1.1450 ;
        RECT  7.2750 0.6400 7.3950 1.3800 ;
        RECT  7.1750 1.2600 7.2950 2.2100 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 7.5400 0.1800 ;
        RECT  6.8550 -0.1800 6.9750 0.6900 ;
        RECT  4.5450 0.3500 4.7850 0.4700 ;
        RECT  4.5450 -0.1800 4.6650 0.4700 ;
        RECT  3.7050 -0.1800 3.8250 0.6400 ;
        RECT  1.5450 -0.1800 1.7850 0.3400 ;
        RECT  0.1400 -0.1800 0.2600 0.7150 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 7.5400 2.7900 ;
        RECT  6.6950 2.0300 6.9350 2.1500 ;
        RECT  6.6950 2.0300 6.8150 2.7900 ;
        RECT  4.3500 2.2700 4.5900 2.7900 ;
        RECT  3.6900 2.2100 3.8100 2.7900 ;
        RECT  1.4250 2.0600 1.5450 2.7900 ;
        RECT  0.1400 1.5550 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.1550 1.1400 6.9750 1.1400 6.9750 1.9100 6.0150 1.9100 6.0150 2.0900 5.8950 2.0900
                 5.8950 1.9100 5.6700 1.9100 5.6700 1.9900 5.4300 1.9900 5.4300 1.8700 5.5500 1.8700
                 5.5500 1.7900 6.8550 1.7900 6.8550 0.9300 6.6150 0.9300 6.6150 0.6300 5.6250 0.6300
                 5.6250 0.6400 5.5050 0.6400 5.5050 0.4000 5.6250 0.4000 5.6250 0.5100 6.7350 0.5100
                 6.7350 0.8100 6.9750 0.8100 6.9750 1.0200 7.1550 1.0200 ;
        POLYGON  5.7700 1.6700 5.3100 1.6700 5.3100 2.1500 4.0500 2.1500 4.0500 2.0900 3.7850 2.0900
                 3.7850 2.0300 2.6500 2.0300 2.6500 1.9600 1.6650 1.9600 1.6650 1.9400 0.8250 1.9400
                 0.8250 1.1950 0.3400 1.1950 0.3400 1.0750 0.8250 1.0750 0.8250 0.5000 2.3850 0.5000
                 2.3850 0.4100 3.1250 0.4100 3.1250 0.4600 3.2450 0.4600 3.2450 0.5800 3.0050 0.5800
                 3.0050 0.5300 2.5050 0.5300 2.5050 0.9200 2.3850 0.9200 2.3850 0.6200 0.9450 0.6200
                 0.9450 1.8200 1.7850 1.8200 1.7850 1.8400 2.3850 1.8400 2.3850 1.6600 2.5050 1.6600
                 2.5050 1.8400 2.7700 1.8400 2.7700 1.9100 2.9900 1.9100 2.9900 1.7900 3.1100 1.7900
                 3.1100 1.9100 3.9050 1.9100 3.9050 1.9700 4.1700 1.9700 4.1700 2.0300 5.1900 2.0300
                 5.1900 1.5500 5.7700 1.5500 ;
        POLYGON  5.2050 0.7100 4.1250 0.7100 4.1250 0.4000 4.2450 0.4000 4.2450 0.5900 5.0850 0.5900
                 5.0850 0.4000 5.2050 0.4000 ;
        POLYGON  5.0700 1.9100 4.8300 1.9100 4.8300 1.8500 4.0500 1.8500 4.0500 1.6100 4.1700 1.6100
                 4.1700 1.7300 4.9500 1.7300 4.9500 1.7900 5.0700 1.7900 ;
        RECT  1.0650 0.7400 2.1450 0.8600 ;
        POLYGON  2.1450 1.7200 1.9050 1.7200 1.9050 1.7000 1.0650 1.7000 1.0650 1.5800 2.0250 1.5800
                 2.0250 1.6000 2.1450 1.6000 ;
    END
END ADDFX1

MACRO ADDFHXL
    CLASS CORE ;
    FOREIGN ADDFHXL 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2580  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.1400 0.8700 6.2350 0.9900 ;
        RECT  4.1400 0.8000 4.2600 1.0600 ;
        RECT  4.1150 0.8700 6.2350 0.9200 ;
        RECT  3.7500 0.7800 4.2350 0.9000 ;
        RECT  2.9350 0.7500 3.8700 0.8700 ;
        RECT  2.9150 0.6500 3.1750 0.8000 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3440  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.9750 1.2300 7.2350 1.3800 ;
        RECT  4.8350 1.1100 7.2150 1.2300 ;
        RECT  5.0650 1.1100 5.1850 1.3500 ;
        RECT  3.6550 1.1800 5.1850 1.3000 ;
        RECT  3.6550 1.0200 3.8950 1.3000 ;
        RECT  3.5100 1.0200 3.8950 1.1400 ;
        RECT  1.6950 0.9900 3.6300 1.1000 ;
        RECT  2.4900 1.0200 3.8950 1.1100 ;
        RECT  1.6950 0.9800 2.6100 1.1000 ;
        RECT  1.6950 0.9800 1.8150 1.2400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3440  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3050 1.3500 6.8550 1.4700 ;
        RECT  4.7750 1.4700 5.4250 1.5900 ;
        RECT  3.3200 1.4200 4.8950 1.5400 ;
        RECT  3.3200 1.2600 3.4850 1.5400 ;
        RECT  2.9150 1.2600 3.4850 1.3800 ;
        RECT  2.0550 1.2400 3.1750 1.3400 ;
        RECT  2.9150 1.2300 3.1750 1.3800 ;
        RECT  2.1750 1.2600 3.4850 1.3600 ;
        RECT  2.0550 1.2200 2.2950 1.3400 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2408  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5600 1.3650 0.6800 2.1250 ;
        RECT  0.0700 0.8850 0.6800 1.0050 ;
        RECT  0.5600 0.6250 0.6800 1.0050 ;
        RECT  0.1000 1.3650 0.6800 1.4850 ;
        RECT  0.1000 0.8850 0.2200 1.4850 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.2408  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.7150 1.4650 8.0500 1.7250 ;
        RECT  7.7150 0.5000 7.8350 2.2100 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.1750 0.3900 7.4150 0.5100 ;
        RECT  7.1750 -0.1800 7.2950 0.5100 ;
        RECT  4.8350 0.3900 5.0750 0.5100 ;
        RECT  4.8350 -0.1800 4.9550 0.5100 ;
        RECT  3.9950 -0.1800 4.1150 0.6400 ;
        RECT  1.7150 -0.1800 1.9550 0.3800 ;
        RECT  0.1400 -0.1800 0.2600 0.7650 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.1750 2.0700 7.4150 2.1900 ;
        RECT  7.1750 2.0700 7.2950 2.7900 ;
        RECT  4.8250 2.2900 5.0650 2.7900 ;
        RECT  3.8650 1.9000 3.9850 2.7900 ;
        RECT  3.7450 1.9000 3.9850 2.1500 ;
        RECT  1.7150 2.2200 1.9550 2.7900 ;
        RECT  0.1400 1.6050 0.2600 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.5950 1.5500 7.4750 1.5500 7.4750 1.9500 6.2950 1.9500 6.2950 2.2100 6.1750 2.2100
                 6.1750 1.9500 5.9050 1.9500 5.9050 2.1700 5.7850 2.1700 5.7850 1.8300 7.3550 1.8300
                 7.3550 0.7500 5.7950 0.7500 5.7950 0.4900 5.9150 0.4900 5.9150 0.6300 6.3150 0.6300
                 6.3150 0.4900 6.4350 0.4900 6.4350 0.6300 7.4750 0.6300 7.4750 1.4300 7.5950 1.4300 ;
        POLYGON  6.0850 1.7100 5.6650 1.7100 5.6650 2.1700 4.1050 2.1700 4.1050 1.7800 3.5500 1.7800
                 3.5500 2.0000 3.2850 2.0000 3.2850 2.2100 3.1650 2.2100 3.1650 2.0000 2.7950 2.0000
                 2.7950 2.1000 0.9950 2.1000 0.9950 1.2450 0.3400 1.2450 0.3400 1.1250 0.9950 1.1250
                 0.9950 0.5000 2.6750 0.5000 2.6750 0.4100 3.4150 0.4100 3.4150 0.4600 3.5350 0.4600
                 3.5350 0.5800 3.2950 0.5800 3.2950 0.5300 2.7950 0.5300 2.7950 0.8200 2.6750 0.8200
                 2.6750 0.6200 1.1150 0.6200 1.1150 1.9800 2.6750 1.9800 2.6750 1.4800 2.7950 1.4800
                 2.7950 1.8800 3.1650 1.8800 3.1650 1.6900 3.2850 1.6900 3.2850 1.8800 3.4300 1.8800
                 3.4300 1.6600 4.2250 1.6600 4.2250 2.0500 5.5450 2.0500 5.5450 1.5900 6.0850 1.5900 ;
        POLYGON  5.4950 0.7500 4.4750 0.7500 4.4750 0.6800 4.3550 0.6800 4.3550 0.5600 4.5950 0.5600
                 4.5950 0.6300 5.3750 0.6300 5.3750 0.5000 5.4950 0.5000 ;
        POLYGON  5.4250 1.8900 5.1850 1.8900 5.1850 1.8600 4.5850 1.8600 4.5850 1.9300 4.3450 1.9300
                 4.3450 1.7400 5.1850 1.7400 5.1850 1.7100 5.4250 1.7100 ;
        RECT  1.2350 0.7400 2.4350 0.8600 ;
        POLYGON  2.3750 1.8600 2.2550 1.8600 2.2550 1.6000 1.5350 1.6000 1.5350 1.8600 1.4150 1.8600
                 1.4150 1.3400 1.5350 1.3400 1.5350 1.4800 2.3750 1.4800 ;
    END
END ADDFHXL

MACRO ADDFHX4
    CLASS CORE ;
    FOREIGN ADDFHX4 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 10.4400 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3240  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.0350 0.8200 7.4950 0.9400 ;
        RECT  5.1750 0.8200 5.4150 1.0900 ;
        RECT  4.0550 0.7800 5.1550 0.9000 ;
        RECT  4.0750 0.6500 4.3350 0.9000 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.2750 0.9400 8.3950 1.2500 ;
        RECT  8.1350 0.9400 8.3950 1.1600 ;
        RECT  7.6550 1.0400 8.3950 1.1600 ;
        RECT  5.5350 1.0600 7.7750 1.1800 ;
        RECT  4.7950 1.2100 5.6550 1.3300 ;
        RECT  5.5350 1.0600 5.6550 1.3300 ;
        RECT  4.7950 1.0200 4.9150 1.3300 ;
        RECT  3.7350 1.0200 4.9150 1.1400 ;
        RECT  2.6750 0.9800 3.8550 1.1000 ;
        RECT  2.6750 0.9800 2.7950 1.2400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.4320  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.8950 1.2800 8.1350 1.4000 ;
        RECT  5.7750 1.3000 8.0150 1.4200 ;
        RECT  4.4200 1.4500 5.8950 1.5700 ;
        RECT  5.7750 1.3000 5.8950 1.5700 ;
        RECT  4.4200 1.2800 4.6750 1.5700 ;
        RECT  4.4200 1.2800 4.5700 1.7250 ;
        RECT  4.0500 1.2800 4.6750 1.4000 ;
        RECT  3.1350 1.2600 4.1700 1.3400 ;
        RECT  3.2550 1.2800 4.6750 1.3800 ;
        RECT  3.1350 1.2200 3.3750 1.3400 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  1.4350 1.3200 1.5550 2.2100 ;
        RECT  1.4350 0.6700 1.5550 0.9600 ;
        RECT  0.5550 1.3200 1.5550 1.4400 ;
        RECT  0.5550 0.8400 1.5550 0.9600 ;
        RECT  0.5950 1.3200 0.7150 2.2100 ;
        RECT  0.5950 0.6700 0.7150 0.9600 ;
        RECT  0.5550 0.7900 0.6750 1.4400 ;
        RECT  0.3600 0.8850 0.6750 1.1450 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.6912  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  9.7350 0.8850 10.0800 1.1450 ;
        RECT  8.8550 1.3200 9.8550 1.4400 ;
        RECT  9.7350 0.7600 9.8550 1.4400 ;
        RECT  9.6950 1.3200 9.8150 2.2100 ;
        RECT  8.8550 0.7600 9.8550 0.8800 ;
        RECT  9.6950 0.5900 9.8150 0.8800 ;
        RECT  8.8550 1.3200 8.9750 2.2100 ;
        RECT  8.8550 0.5900 8.9750 0.8800 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 10.4400 0.1800 ;
        RECT  10.1150 -0.1800 10.2350 0.6400 ;
        RECT  9.2750 -0.1800 9.3950 0.6400 ;
        RECT  8.3750 0.4600 8.6150 0.5800 ;
        RECT  8.3750 -0.1800 8.4950 0.5800 ;
        RECT  5.9350 0.3400 6.1750 0.4600 ;
        RECT  5.9350 -0.1800 6.0550 0.4600 ;
        RECT  5.0950 -0.1800 5.2150 0.6400 ;
        RECT  2.8150 -0.1800 3.0550 0.3800 ;
        RECT  1.8550 -0.1800 1.9750 0.7200 ;
        RECT  1.0150 -0.1800 1.1350 0.7200 ;
        RECT  0.1750 -0.1800 0.2950 0.7200 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 10.4400 2.7900 ;
        RECT  10.1150 1.5600 10.2350 2.7900 ;
        RECT  9.2750 1.5600 9.3950 2.7900 ;
        RECT  8.3750 2.0200 8.6150 2.1500 ;
        RECT  8.3750 2.0200 8.4950 2.7900 ;
        RECT  5.9350 2.1700 6.1750 2.7900 ;
        RECT  4.9750 2.1700 5.2150 2.7900 ;
        RECT  2.8750 2.1000 2.9950 2.7900 ;
        RECT  1.7950 2.0300 2.0350 2.1500 ;
        RECT  1.7950 2.0300 1.9150 2.7900 ;
        RECT  1.0150 1.5600 1.1350 2.7900 ;
        RECT  0.1750 1.5600 0.2950 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  9.6150 1.1200 8.6350 1.1200 8.6350 1.9000 7.6550 1.9000 7.6550 2.1500 7.4150 2.1500
                 7.4150 1.9000 7.2550 1.9000 7.2550 2.1500 7.0150 2.1500 7.0150 1.8800 7.1350 1.8800
                 7.1350 1.7800 8.5150 1.7800 8.5150 0.8200 8.1350 0.8200 8.1350 0.7000 6.8350 0.7000
                 6.8350 0.5800 7.5150 0.5800 7.5150 0.5000 7.7550 0.5000 7.7550 0.5800 8.2550 0.5800
                 8.2550 0.7000 8.6350 0.7000 8.6350 1.0000 9.6150 1.0000 ;
        POLYGON  7.3350 1.6600 6.8950 1.6600 6.8950 2.0500 4.4550 2.0500 4.4550 2.2100 4.3350 2.2100
                 4.3350 2.0500 3.8950 2.0500 3.8950 2.1500 3.7750 2.1500 3.7750 2.0500 3.6850 2.0500
                 3.6850 1.9800 2.3600 1.9800 2.3600 1.9100 2.0950 1.9100 2.0950 1.2000 0.7950 1.2000
                 0.7950 1.0800 2.0950 1.0800 2.0950 0.5000 3.7750 0.5000 3.7750 0.4100 4.5750 0.4100
                 4.5750 0.6500 4.4550 0.6500 4.4550 0.5300 3.8950 0.5300 3.8950 0.7400 3.7750 0.7400
                 3.7750 0.6200 2.2150 0.6200 2.2150 1.7900 2.4800 1.7900 2.4800 1.8600 3.7750 1.8600
                 3.7750 1.5000 3.8950 1.5000 3.8950 1.9300 4.3350 1.9300 4.3350 1.8450 4.4550 1.8450
                 4.4550 1.9300 6.7750 1.9300 6.7750 1.5400 7.3350 1.5400 ;
        RECT  5.4550 0.5800 6.6550 0.7000 ;
        POLYGON  6.6550 1.8100 5.4550 1.8100 5.4550 1.6900 6.4150 1.6900 6.4150 1.6200 6.6550 1.6200 ;
        RECT  2.3350 0.7400 3.5350 0.8600 ;
        POLYGON  3.4750 1.7400 3.3550 1.7400 3.3550 1.6200 2.5150 1.6200 2.5150 1.6700 2.3950 1.6700
                 2.3950 1.3400 2.5150 1.3400 2.5150 1.5000 3.4750 1.5000 ;
    END
END ADDFHX4

MACRO ADDFHX2
    CLASS CORE ;
    FOREIGN ADDFHX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.7000 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2580  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.5050 0.8300 6.5450 0.9500 ;
        RECT  4.5650 0.8200 4.6850 1.0600 ;
        RECT  3.2050 0.7800 3.6250 0.9000 ;
        RECT  3.2050 0.6500 3.4650 0.9000 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3440  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.3250 1.0700 7.4450 1.3100 ;
        RECT  5.0950 1.0700 7.4450 1.1900 ;
        RECT  6.9750 0.9400 7.2350 1.1900 ;
        RECT  4.3250 1.1800 5.2150 1.3000 ;
        RECT  3.0650 1.0700 4.4450 1.1900 ;
        RECT  2.8000 1.0200 3.1850 1.1400 ;
        RECT  2.0050 0.9900 2.9200 1.1100 ;
        RECT  1.8850 1.0600 2.1250 1.1800 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3440  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  5.3350 1.3100 7.1650 1.4300 ;
        RECT  2.9150 1.4200 5.4550 1.5400 ;
        RECT  2.9150 1.3100 3.1750 1.6700 ;
        RECT  2.7900 1.3100 3.1750 1.4300 ;
        RECT  2.2850 1.2600 2.9100 1.3500 ;
        RECT  2.5250 1.3100 3.1750 1.3800 ;
        RECT  2.2850 1.2300 2.6450 1.3500 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5850 0.6800 0.7050 2.2100 ;
        RECT  0.3600 0.8850 0.7050 1.1450 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3456  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  8.0250 0.8850 8.3400 1.1450 ;
        RECT  8.0250 0.5900 8.1450 1.6800 ;
        RECT  7.9050 1.5600 8.0250 2.2100 ;
        END
    END S
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.7000 0.1800 ;
        RECT  8.4450 -0.1800 8.5650 0.6400 ;
        RECT  7.4850 0.3500 7.7250 0.4700 ;
        RECT  7.4850 -0.1800 7.6050 0.4700 ;
        RECT  5.0650 0.3500 5.3050 0.4700 ;
        RECT  5.0650 -0.1800 5.1850 0.4700 ;
        RECT  4.2250 -0.1800 4.3450 0.6400 ;
        RECT  1.9650 -0.1800 2.2050 0.3800 ;
        RECT  1.0050 -0.1800 1.1250 0.7300 ;
        RECT  0.1650 -0.1800 0.2850 0.7300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.7000 2.7900 ;
        RECT  8.3250 1.5600 8.4450 2.7900 ;
        RECT  7.4250 2.0300 7.6650 2.1500 ;
        RECT  7.4250 2.0300 7.5450 2.7900 ;
        RECT  5.2250 2.2300 5.3450 2.7900 ;
        RECT  4.2050 2.2200 4.4450 2.7900 ;
        RECT  1.9650 2.2000 2.2050 2.7900 ;
        RECT  1.0650 1.9800 1.1850 2.7900 ;
        RECT  0.1650 1.5600 0.2850 2.7900 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        POLYGON  7.8850 1.4400 7.6850 1.4400 7.6850 1.9100 6.6050 1.9100 6.6050 2.2100 6.4850 2.2100
                 6.4850 1.9100 6.1850 1.9100 6.1850 2.0700 6.0650 2.0700 6.0650 1.7900 7.5650 1.7900
                 7.5650 0.7100 6.0850 0.7100 6.0850 0.6300 5.9650 0.6300 5.9650 0.5100 6.2050 0.5100
                 6.2050 0.5900 6.6250 0.5900 6.6250 0.4500 6.7450 0.4500 6.7450 0.5900 7.6850 0.5900
                 7.6850 1.2000 7.8850 1.2000 ;
        POLYGON  6.4250 1.6700 5.9450 1.6700 5.9450 2.1100 4.8900 2.1100 4.8900 2.1000 3.6850 2.1000
                 3.6850 2.2000 3.5650 2.2000 3.5650 2.1000 2.9250 2.1000 2.9250 2.0800 1.5100 2.0800
                 1.5100 1.8600 1.2450 1.8600 1.2450 1.2600 0.8250 1.2600 0.8250 1.1400 1.2450 1.1400
                 1.2450 0.5000 2.9250 0.5000 2.9250 0.4100 3.5850 0.4100 3.5850 0.4000 3.7050 0.4000
                 3.7050 0.6400 3.5850 0.6400 3.5850 0.5300 3.0450 0.5300 3.0450 0.8200 2.9250 0.8200
                 2.9250 0.6200 1.3650 0.6200 1.3650 1.7400 1.6300 1.7400 1.6300 1.9600 2.9250 1.9600
                 2.9250 1.7900 3.0450 1.7900 3.0450 1.9800 3.5650 1.9800 3.5650 1.6800 3.6850 1.6800
                 3.6850 1.9800 5.0100 1.9800 5.0100 1.9900 5.8250 1.9900 5.8250 1.5500 6.4250 1.5500 ;
        POLYGON  5.7250 0.7100 4.8050 0.7100 4.8050 0.6800 4.5850 0.6800 4.5850 0.5600 4.9250 0.5600
                 4.9250 0.5900 5.6050 0.5900 5.6050 0.4700 5.7250 0.4700 ;
        POLYGON  5.7050 1.8700 5.5850 1.8700 5.5850 1.8600 4.6850 1.8600 4.6850 1.7400 5.5850 1.7400
                 5.5850 1.5500 5.7050 1.5500 ;
        RECT  1.4850 0.7400 2.6850 0.8600 ;
        POLYGON  2.6850 1.8400 2.4450 1.8400 2.4450 1.6200 1.6650 1.6200 1.6650 1.3400 1.7850 1.3400
                 1.7850 1.5000 2.5650 1.5000 2.5650 1.5700 2.6850 1.5700 ;
    END
END ADDFHX2

MACRO ADDFHX1
    CLASS CORE ;
    FOREIGN ADDFHX1 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.1200 BY 2.6100 ;
    SYMMETRY X Y ;
    SITE gsclib090site ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  7.5850 0.8850 7.7600 1.1450 ;
        RECT  7.5850 0.5900 7.7050 2.2100 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.3024  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.5600 1.3200 0.6800 2.2100 ;
        RECT  0.5600 0.6700 0.6800 0.9600 ;
        RECT  0.1000 1.3200 0.6800 1.4400 ;
        RECT  0.1000 0.8400 0.6800 0.9600 ;
        RECT  0.1000 0.8400 0.2200 1.4400 ;
        RECT  0.0700 0.8850 0.2200 1.1450 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3440  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.5000 1.3700 6.6200 1.6100 ;
        RECT  4.7450 1.3900 6.6200 1.5100 ;
        RECT  3.1600 1.4400 4.8650 1.5400 ;
        RECT  4.3600 1.4200 6.6200 1.5100 ;
        RECT  3.1600 1.4400 4.6000 1.5600 ;
        RECT  3.1600 1.2800 3.4000 1.5600 ;
        RECT  1.9900 1.2200 3.2800 1.3400 ;
        RECT  2.9150 1.2800 3.4000 1.3800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.3440  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  6.7700 1.1100 7.0850 1.2300 ;
        RECT  6.7400 1.1300 6.8900 1.4350 ;
        RECT  6.2600 1.1300 6.8900 1.2500 ;
        RECT  3.5900 1.1800 6.3800 1.2700 ;
        RECT  4.5050 1.1500 7.0850 1.2300 ;
        RECT  3.5900 1.1800 4.6250 1.3000 ;
        RECT  3.5900 1.0200 3.8300 1.3200 ;
        RECT  3.4450 1.0200 3.8300 1.1400 ;
        RECT  1.5900 0.9800 3.5650 1.1000 ;
        RECT  1.4700 1.0600 1.7100 1.1800 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.2580  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  4.0750 0.9100 6.1400 1.0300 ;
        RECT  4.0750 0.7800 4.1950 1.0600 ;
        RECT  3.6850 0.7800 4.1950 0.9000 ;
        RECT  2.8900 0.7400 3.8050 0.8600 ;
        RECT  2.9150 0.6500 3.1750 0.8600 ;
        END
    END CI
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 8.1200 2.7900 ;
        RECT  7.0450 2.1100 7.2850 2.2300 ;
        RECT  7.0450 2.1100 7.1650 2.7900 ;
        RECT  4.7400 2.2300 4.8600 2.7900 ;
        RECT  3.7200 2.2200 3.9600 2.7900 ;
        RECT  1.6700 1.9400 1.9100 2.7900 ;
        RECT  0.1400 1.5600 0.2600 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 8.1200 0.1800 ;
        RECT  7.0450 0.4300 7.2850 0.5500 ;
        RECT  7.0450 -0.1800 7.1650 0.5500 ;
        RECT  4.8350 0.4300 5.0750 0.5500 ;
        RECT  4.8350 -0.1800 4.9550 0.5500 ;
        RECT  3.9950 -0.1800 4.1150 0.6400 ;
        RECT  1.6700 -0.1800 1.9100 0.3800 ;
        RECT  0.1400 -0.1800 0.2600 0.7200 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  7.4650 1.3850 7.3250 1.3850 7.3250 1.9900 6.1200 1.9900 6.1200 2.2100 6.0000 2.2100
                 6.0000 1.9900 5.7000 1.9900 5.7000 2.1500 5.5800 2.1500 5.5800 1.8700 7.2050 1.8700
                 7.2050 0.7900 5.8550 0.7900 5.8550 0.6800 5.7350 0.6800 5.7350 0.5600 5.9750 0.5600
                 5.9750 0.6700 6.1850 0.6700 6.1850 0.5000 6.3050 0.5000 6.3050 0.6700 7.3250 0.6700
                 7.3250 1.2650 7.4650 1.2650 ;
        POLYGON  5.9400 1.7500 5.4600 1.7500 5.4600 2.1100 4.6700 2.1100 4.6700 2.1000 3.2000 2.1000
                 3.2000 2.2000 3.0800 2.2000 3.0800 2.1000 2.6300 2.1000 2.6300 2.2500 2.0300 2.2500
                 2.0300 1.8200 0.9500 1.8200 0.9500 1.2000 0.3400 1.2000 0.3400 1.0800 0.9500 1.0800
                 0.9500 0.5000 2.6300 0.5000 2.6300 0.4100 3.4150 0.4100 3.4150 0.4600 3.5350 0.4600
                 3.5350 0.5800 3.2950 0.5800 3.2950 0.5300 2.7500 0.5300 2.7500 0.8200 2.6300 0.8200
                 2.6300 0.6200 1.0700 0.6200 1.0700 1.7000 2.1500 1.7000 2.1500 2.1300 2.5100 2.1300
                 2.5100 1.9800 2.6900 1.9800 2.6900 1.5000 2.8100 1.5000 2.8100 1.9800 3.0800 1.9800
                 3.0800 1.6800 3.2000 1.6800 3.2000 1.9800 4.7900 1.9800 4.7900 1.9900 5.3400 1.9900
                 5.3400 1.6300 5.9400 1.6300 ;
        POLYGON  5.4950 0.7900 4.4750 0.7900 4.4750 0.6800 4.3550 0.6800 4.3550 0.5600 4.5950 0.5600
                 4.5950 0.6700 5.3750 0.6700 5.3750 0.5000 5.4950 0.5000 ;
        POLYGON  5.2200 1.8700 5.1000 1.8700 5.1000 1.8600 4.2000 1.8600 4.2000 1.7400 5.1000 1.7400
                 5.1000 1.6300 5.2200 1.6300 ;
        RECT  1.1900 0.7400 2.3900 0.8600 ;
        POLYGON  2.3900 2.0100 2.2700 2.0100 2.2700 1.5800 1.2500 1.5800 1.2500 1.3400 1.3700 1.3400
                 1.3700 1.4600 2.3900 1.4600 ;
    END
END ADDFHX1

MACRO ACHCONX2
    CLASS CORE ;
    FOREIGN ACHCONX2 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 14.5000 BY 2.6100 ;
    SYMMETRY X Y R90 ;
    SITE gsclib090site ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1940  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  13.5400 1.0800 14.0600 1.3200 ;
        RECT  13.6450 1.0800 13.9050 1.3800 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.7841  LAYER Metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.7200  LAYER Metal1  ;
        ANTENNAMAXAREACAR 1.0890  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  3.1650 1.1300 3.5100 1.4900 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.1940  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  0.1900 1.2300 0.5650 1.3800 ;
        RECT  0.1900 0.9750 0.4300 1.3800 ;
        END
    END A
    PIN CON
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.1716  LAYER Metal1  ;
        PORT
        LAYER Metal1 ;
        RECT  11.9700 1.5700 12.9300 1.6900 ;
        RECT  10.5300 0.3600 12.9300 0.4800 ;
        RECT  11.9050 1.2300 12.1650 1.3800 ;
        RECT  10.5300 1.8050 12.0900 1.9250 ;
        RECT  11.9700 0.3600 12.0900 1.9250 ;
        END
    END CON
    PIN VDD
        DIRECTION INPUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 2.4300 14.5000 2.7900 ;
        RECT  14.1600 1.7100 14.4000 2.7900 ;
        RECT  13.0800 2.1400 13.3200 2.7900 ;
        RECT  10.1400 2.2900 10.3800 2.7900 ;
        RECT  9.0600 2.2900 9.3000 2.7900 ;
        RECT  3.3300 2.2900 3.5700 2.7900 ;
        RECT  2.2500 2.2900 2.4900 2.7900 ;
        RECT  1.1700 1.7100 1.4100 2.7900 ;
        RECT  0.0900 1.7700 0.3300 2.7900 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  0.0000 -0.1800 14.5000 0.1800 ;
        RECT  14.1600 -0.1800 14.4000 0.7250 ;
        RECT  13.0800 -0.1800 13.3200 0.5800 ;
        RECT  10.1400 -0.1800 10.3800 0.3200 ;
        RECT  9.0600 -0.1800 9.3000 0.3200 ;
        RECT  3.3300 -0.1800 3.5700 0.3200 ;
        RECT  2.2500 -0.1800 2.4900 0.3200 ;
        RECT  1.1700 -0.1800 1.4100 0.6400 ;
        RECT  0.0900 -0.1800 0.3300 0.6400 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        POLYGON  13.8600 0.5600 13.7400 0.5600 13.7400 0.8600 13.1700 0.8600 13.1700 1.6550
                 13.8600 1.6550 13.8600 2.1500 13.6200 2.1500 13.6200 1.7750 13.1700 1.7750
                 13.1700 1.9300 12.3900 1.9300 12.3900 2.2500 12.1500 2.2500 12.1500 2.1300
                 12.2100 2.1300 12.2100 1.8100 13.0500 1.8100 13.0500 0.8600 12.3900 0.8600
                 12.3900 0.9200 12.2100 0.9200 12.2100 0.6800 12.3900 0.6800 12.3900 0.7400
                 13.6200 0.7400 13.6200 0.4400 13.8600 0.4400 ;
        POLYGON  11.8500 1.0950 11.6600 1.0950 11.6600 1.3300 11.0000 1.3300 11.0000 1.4100
                 10.8800 1.4100 10.8800 1.6850 10.4100 1.6850 10.4100 1.9300 9.3300 1.9300
                 9.3300 1.7700 6.4800 1.7700 6.4800 1.5300 5.3400 1.5300 5.3400 1.4100 5.4300 1.4100
                 5.4300 0.7200 5.3400 0.7200 5.3400 0.6000 7.0500 0.6000 7.0500 0.7200 5.5500 0.7200
                 5.5500 1.4100 6.6000 1.4100 6.6000 1.6500 9.4500 1.6500 9.4500 1.8100 10.2900 1.8100
                 10.2900 1.5650 10.7600 1.5650 10.7600 1.2100 11.5400 1.2100 11.5400 0.7850
                 11.8500 0.7850 ;
        POLYGON  11.3100 0.7200 10.6400 0.7200 10.6400 1.2800 9.8400 1.2800 9.8400 1.6900 9.6000 1.6900
                 9.6000 1.5700 9.7200 1.5700 9.7200 0.8600 9.6000 0.8600 9.6000 0.7400 9.8400 0.7400
                 9.8400 1.1600 10.5200 1.1600 10.5200 0.6000 11.3100 0.6000 ;
        POLYGON  11.3100 2.1700 9.8400 2.1700 9.8400 2.2500 9.6000 2.2500 9.6000 2.0500 11.3100 2.0500 ;
        POLYGON  10.4000 0.9850 10.1600 0.9850 10.1600 0.5600 9.4800 0.5600 9.4800 0.7200 8.3100 0.7200
                 8.3100 1.4100 8.3700 1.4100 8.3700 1.5300 8.1300 1.5300 8.1300 1.4100 8.1900 1.4100
                 8.1900 0.7200 8.1300 0.7200 8.1300 0.6000 9.3600 0.6000 9.3600 0.4400 10.2800 0.4400
                 10.2800 0.8650 10.4000 0.8650 ;
        POLYGON  9.4150 1.4250 8.8750 1.4250 8.8750 0.9850 8.6550 0.9850 8.6550 0.8650 8.9950 0.8650
                 8.9950 1.3050 9.1650 1.3050 9.1650 0.9850 9.4150 0.9850 ;
        POLYGON  8.9100 0.4800 8.0100 0.4800 8.0100 1.5300 7.3700 1.5300 7.3700 1.4100 7.8900 1.4100
                 7.8900 0.4800 6.2700 0.4800 6.2700 0.3600 8.9100 0.3600 ;
        POLYGON  8.9100 2.2500 3.6900 2.2500 3.6900 2.1700 2.1350 2.1700 2.1350 2.2500 1.7100 2.2500
                 1.7100 2.1300 1.7700 2.1300 1.7700 0.6850 1.7100 0.6850 1.7100 0.5650 1.9500 0.5650
                 1.9500 0.6850 1.8900 0.6850 1.8900 2.1300 2.0150 2.1300 2.0150 2.0500 3.8100 2.0500
                 3.8100 2.1300 8.9100 2.1300 ;
        POLYGON  8.3700 2.0100 6.2400 2.0100 6.2400 1.7700 4.1650 1.7700 4.1650 1.6850 4.0000 1.6850
                 4.0000 1.0500 4.0800 1.0500 4.0800 0.6000 4.5000 0.6000 4.5000 0.7200 4.2000 0.7200
                 4.2000 1.1700 4.1200 1.1700 4.1200 1.5650 4.2850 1.5650 4.2850 1.6500 6.3600 1.6500
                 6.3600 1.8900 8.3700 1.8900 ;
        POLYGON  7.7700 1.2900 7.5500 1.2900 7.5500 1.1250 6.9800 1.1250 6.9800 0.9600 6.3250 0.9600
                 6.3250 0.8400 7.1000 0.8400 7.1000 1.0050 7.7700 1.0050 ;
        POLYGON  7.0300 1.4900 6.7900 1.4900 6.7900 1.3650 6.7150 1.3650 6.7150 1.2900 5.8000 1.2900
                 5.8000 1.0250 5.6800 1.0250 5.6800 0.8400 5.9200 0.8400 5.9200 1.1700 6.8350 1.1700
                 6.8350 1.2450 7.0300 1.2450 ;
        POLYGON  6.1200 0.4800 3.9600 0.4800 3.9600 0.5600 2.3850 0.5600 2.3850 1.8100 4.0450 1.8100
                 4.0450 1.8900 6.1200 1.8900 6.1200 2.0100 3.9250 2.0100 3.9250 1.9300 2.2650 1.9300
                 2.2650 1.2500 2.0500 1.2500 2.0500 1.1300 2.2650 1.1300 2.2650 0.4400 3.7200 0.4400
                 3.7200 0.3600 6.1200 0.3600 ;
        POLYGON  5.0800 1.4250 4.2400 1.4250 4.2400 1.3050 4.9600 1.3050 4.9600 1.0250 4.9000 1.0250
                 4.9000 0.7300 5.0800 0.7300 ;
        POLYGON  3.8800 0.9850 3.6400 0.9850 3.6400 0.8750 2.9700 0.8750 2.9700 1.5700 3.0300 1.5700
                 3.0300 1.6900 2.7900 1.6900 2.7900 1.5700 2.8500 1.5700 2.8500 0.8750 2.7900 0.8750
                 2.7900 0.7400 3.0300 0.7400 3.0300 0.7550 3.8800 0.7550 ;
        POLYGON  1.5100 1.2500 0.8100 1.2500 0.8100 1.6250 0.8700 1.6250 0.8700 2.0650 0.6300 2.0650
                 0.6300 1.6250 0.6900 1.6250 0.6900 0.6850 0.6300 0.6850 0.6300 0.5650 0.8700 0.5650
                 0.8700 0.6850 0.8100 0.6850 0.8100 1.1300 1.5100 1.1300 ;
    END
END ACHCONX2

END LIBRARY
