# Important Info: This tech-Lef file define vias (but not metal layers which already 
#                 defined from "gpdk090" techlib.)
#
#
# NOTE!!!  These statements are ORDER DEPENDENT.  Refer to LEF syntax documentation.
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

# "LEF" format is always in microns (DEF uses this).
UNITS 
  #DATABASE MICRONS 100 ; # Soc-E default
  DATABASE MICRONS 2000 ;
#  CAPACITANCE PICOFARADS 1 ;#Commented out since it is already specified in gpdk090_oa.tf
END UNITS
#
#
SITE gsclib090site
     SYMMETRY Y  ;
     CLASS core  ;
     SIZE 0.2900 BY 2.6100 ;
END gsclib090site
#


VIA VIA1X DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal1 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal2 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA1X

# Via 2 - for Metal2 pin access (vertical metals)
VIA VIA1V DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal1 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal2 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA1V

# Via 3 - for Metal2 pin access (horizontal metals)
VIA VIA1H DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal1 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal2 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA1H

# Via 4 - for Metal2 pin access (cross rotate)
VIA VIA1XR90 DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal1 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal2 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA1XR90


# Via 5 - double cut east
VIA VIA1_2CUT_E DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal1 ;
    RECT -0.130 -0.075 0.420 0.075 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT  0.220 -0.070 0.360 0.070 ;
  LAYER Metal2 ;
    RECT -0.130 -0.075 0.420 0.075 ;
END VIA1_2CUT_E

# Via 6 - double cut west
VIA VIA1_2CUT_W DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal1 ;
    RECT -0.420 -0.075  0.130 0.075 ;
  LAYER Via1 ;
    RECT -0.360 -0.070 -0.220 0.070 ;
    RECT -0.070 -0.070  0.070 0.070 ;
  LAYER Metal2 ;
    RECT -0.420 -0.075  0.130 0.075 ;
END VIA1_2CUT_W

# Via 7 - double cut north
VIA VIA1_2CUT_N DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal1 ;
    RECT -0.075 -0.130 0.075 0.420 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT -0.070  0.220 0.070 0.360 ;
  LAYER Metal2 ;
    RECT -0.075 -0.130 0.075 0.420 ;
END VIA1_2CUT_N

# Via 8 - double cut south
VIA VIA1_2CUT_S DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal1 ;
    RECT -0.075 -0.420 0.075  0.130 ;
  LAYER Via1 ;
    RECT -0.070 -0.360 0.070 -0.220 ;
    RECT -0.070 -0.070 0.070  0.070 ;
  LAYER Metal2 ;
    RECT -0.075 -0.420 0.075  0.130 ;
END VIA1_2CUT_S

# Via 9 - quad cut square
VIA VIA1_2X2CUT DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal1 ;
    RECT -0.275 -0.220  0.275  0.220 ;
  LAYER Via1 ;
    RECT  0.075  0.075  0.215  0.215 ;
    RECT -0.215  0.075 -0.075  0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT  0.075 -0.215  0.215 -0.075 ;
  LAYER Metal2 ;
    RECT -0.220 -0.275  0.220  0.275 ; 
END VIA1_2X2CUT


# Via 1 - Pin access Metal2 or Metal3
VIA VIA2X DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA2X

# Via 2 - Pin access Metal2 or Metal3
VIA VIA2H DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA2H

# Via 3 - Pin access Metal2 or Metal3
VIA VIA2V DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal3 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA2V

# Via 4 - Pin access Metal2 or Metal3
VIA VIA2XR90 DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal3 ; 
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA2XR90

## Via 5 - TOS via for 3 signal wire
#VIA VIA2TOS DEFAULT
#  TOPOFSTACKONLY
#  RESISTANCE 1.4 ;
#  LAYER Metal2 ;
#    RECT -0.135 -0.170 0.135 0.170 ;
#  LAYER Via2 ;
#    RECT -0.070 -0.070 0.070 0.070 ;
#  LAYER Metal3 ;
#    RECT -0.130 -0.075 0.130 0.075 ;
#END VIA2TOS

VIA VIA2TOS DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.075 -0.27 0.075 0.27 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA2TOS

VIA VIA2TOS_S DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.075 -0.41 0.075 0.13 ;
  LAYER Via2 ;
    RECT -0.070 -0.07 0.070 0.07 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA2TOS_S

VIA VIA2TOS_N DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.41 ;
  LAYER Via2 ;
    RECT -0.070 -0.07 0.070 0.07 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA2TOS_N


# Via 6 - double cut north
VIA VIA2_2CUT_N DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal2 ;
    RECT -0.075 -0.130 0.075 0.420 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT -0.070  0.220 0.070 0.360 ;
  LAYER Metal3 ;
    RECT -0.075 -0.130 0.075 0.420 ;
END VIA2_2CUT_N

# Via 7 - double cut south
VIA VIA2_2CUT_S DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal2 ;
    RECT -0.075 -0.420 0.075  0.130 ;
  LAYER Via2 ;
    RECT -0.070 -0.360 0.070 -0.220 ;
    RECT -0.070 -0.070 0.070  0.070 ;
  LAYER Metal3 ;
    RECT -0.075 -0.420 0.075  0.130 ;
END VIA2_2CUT_S

# Via 8 - double cut east
VIA VIA2_2CUT_E DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal2 ;
    RECT -0.130 -0.075 0.420 0.075 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT  0.220 -0.070 0.360 0.070 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.420 0.075 ;
END VIA2_2CUT_E

# Via 9 - double cut west
VIA VIA2_2CUT_W DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal2 ;
    RECT -0.420 -0.075  0.130 0.075 ;
  LAYER Via2 ;
    RECT -0.360 -0.070 -0.220 0.070 ;
    RECT -0.070 -0.070  0.070 0.070 ;
  LAYER Metal3 ;
    RECT -0.420 -0.075  0.130 0.075 ;
END VIA2_2CUT_W

# Via 10 - quad cut square
VIA VIA2_2X2CUT DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal2 ;     
    RECT -0.220 -0.275  0.220  0.275 ;
  LAYER Via2 ;
    RECT  0.075  0.075  0.215  0.215 ;
    RECT -0.215  0.075 -0.075  0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT  0.075 -0.215  0.215 -0.075 ;
  LAYER Metal3 ;
    RECT -0.275 -0.220  0.275  0.220 ;
END VIA2_2X2CUT


# Via 1 - Pin access Metal3 or Metal4
VIA VIA3X DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA3X

# Via 2 - Pin access Metal3 or Metal4
VIA VIA3H DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA3H

# Via 3 - Pin access Metal3 or Metal4
VIA VIA3V DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA3V

# Via 4 - for Metal3/4 pin access (cross rotate)
VIA VIA3XR90 DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA3XR90


# Via 5 - TOS east no pin access
VIA VIA3TOS_E DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.410 0.075 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA3TOS_E

# Via 6 - TOS west no pin access
VIA VIA3TOS_W DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.410 -0.075 0.130 0.075 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA3TOS_W

# Via 7 - TOS centered no pin access
VIA VIA3TOS DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal3 ;
    RECT -0.270 -0.075 0.270 0.075 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA3TOS

# Via 8 - double cut east
VIA VIA3_2CUT_E DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal3 ;
    RECT -0.130 -0.075 0.420 0.075 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT  0.220 -0.070 0.360 0.070 ;
  LAYER Metal4 ;
    RECT -0.130 -0.075 0.420 0.075 ;
END VIA3_2CUT_E

# Via 9 - double cut west
VIA VIA3_2CUT_W DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal3 ;
    RECT -0.420 -0.075  0.130 0.075 ;
  LAYER Via3 ;
    RECT -0.360 -0.070 -0.220 0.070 ;
    RECT -0.070 -0.070  0.070  0.070 ;
  LAYER Metal4 ;
    RECT -0.420 -0.075  0.130 0.075 ;
END VIA3_2CUT_W

# Via 10 - double cut north
VIA VIA3_2CUT_N DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal3 ;
    RECT -0.075 -0.130 0.075 0.420 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT -0.070  0.220 0.070 0.360 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.420 ;
END VIA3_2CUT_N

# Via 11 - double cut south
VIA VIA3_2CUT_S DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal3 ;
    RECT -0.075 -0.420 0.075  0.130 ;
  LAYER Via3 ;
    RECT -0.070 -0.360 0.070 -0.220 ;
    RECT -0.070 -0.070 0.070  0.070 ;
  LAYER Metal4 ;
    RECT -0.075 -0.420 0.075  0.130 ;
END VIA3_2CUT_S

# Via 12 - quad cut square
VIA VIA3_2X2CUT DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal3 ;
    RECT -0.275 -0.220  0.275  0.220 ;
  LAYER Via3 ;
    RECT  0.075  0.075  0.215  0.215 ;
    RECT -0.215  0.075 -0.075  0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT  0.075 -0.215  0.215 -0.075 ;
  LAYER Metal4 ;
    RECT -0.220 -0.275  0.220  0.275 ;
END VIA3_2X2CUT


# Via 1 - Pin access Metal4 or Metal5
VIA VIA4X DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA4X

# Via 2 - Pin access Metal4 or Metal5
VIA VIA4H DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA4H

# Via 3 - Pin access Metal4 or Metal5
VIA VIA4V DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal5 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA4V

# Via 4 - Pin access Metal4 or Metal5
VIA VIA4XR90 DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal5 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA4XR90

## Via 5 - TOS via for 5 signal wire (no pin access)
#VIA VIA4TOS DEFAULT
#  TOPOFSTACKONLY
#  RESISTANCE 1.4 ;
#  LAYER Metal4 ;
#    RECT -0.135 -0.170 0.135 0.170 ;
#  LAYER Via4 ;
#    RECT -0.070 -0.070 0.070 0.070 ;
#  LAYER Metal5 ;
#    RECT -0.130 -0.075 0.130 0.075 ;
#END VIA4TOS

VIA VIA4TOS DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.075 -0.27 0.075 0.27 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA4TOS

VIA VIA4TOS_S DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.075 -0.41 0.075 0.13 ;
  LAYER Via4 ;
    RECT -0.070 -0.07 0.070 0.07 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA4TOS_S

VIA VIA4TOS_N DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.41 ;
  LAYER Via4 ;
    RECT -0.070 -0.07 0.070 0.07 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA4TOS_N

# Via 6 - double cut north
VIA VIA4_2CUT_N DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal4 ;
    RECT -0.075 -0.130 0.075 0.420 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT -0.070  0.220 0.070 0.360 ;
  LAYER Metal5 ;
    RECT -0.075 -0.130 0.075 0.420 ;
END VIA4_2CUT_N

# Via 7 - double cut south
VIA VIA4_2CUT_S DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal4 ;
    RECT -0.075 -0.420 0.075  0.130 ;
  LAYER Via4 ;
    RECT -0.070 -0.360 0.070 -0.220 ;
    RECT -0.070 -0.070 0.070  0.070 ;
  LAYER Metal5 ;
    RECT -0.075 -0.420 0.075  0.130 ;
END VIA4_2CUT_S

# Via 8 - double cut east
VIA VIA4_2CUT_E DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal4 ;
    RECT -0.130 -0.075 0.420 0.075 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT  0.220 -0.070 0.360 0.070 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.420 0.075 ;
END VIA4_2CUT_E

# Via 9 - double cut west
VIA VIA4_2CUT_W DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal4 ;
    RECT -0.420 -0.075  0.130 0.075 ;
  LAYER Via4 ;
    RECT -0.360 -0.070 -0.220 0.070 ;
    RECT -0.070 -0.070  0.070  0.070 ;
  LAYER Metal5 ;
    RECT -0.420 -0.075  0.130 0.075 ;
END VIA4_2CUT_W

# Via 10 - quad cut square
VIA VIA4_2X2CUT DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal4 ;
    RECT -0.220 -0.275  0.220  0.275 ;
  LAYER Via4 ;
    RECT  0.075  0.075  0.215  0.215 ;
    RECT -0.215  0.075 -0.075  0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT  0.075 -0.215  0.215 -0.075 ;
  LAYER Metal5 ;
    RECT -0.275 -0.220  0.275  0.220 ;
END VIA4_2X2CUT


# Via 1 - Pin access Metal3 or Metal4
VIA VIA5X DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA5X

# Via 2 - Pin access Metal3 or Metal4
VIA VIA5H DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA5H

# Via 3 - Pin access Metal3 or Metal4
VIA VIA5V DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA5V

# Via 4 - for Metal5/6 pin access (cross rotate)
VIA VIA5XR90 DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA5XR90

# Via 5 - TOS east no pin access
VIA VIA5TOS_E DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.410 0.075 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA5TOS_E

# Via 6 - TOS west no pin access
VIA VIA5TOS_W DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.410 -0.075 0.130 0.075 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA5TOS_W

# Via 7 - TOS centered no pin access
VIA VIA5TOS DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal5 ;
    RECT -0.270 -0.075 0.270 0.075 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA5TOS

# Via 8 - double cut east
VIA VIA5_2CUT_E DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal5 ;
    RECT -0.130 -0.075 0.420 0.075 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT  0.220 -0.070 0.360 0.070 ;
  LAYER Metal6 ;
    RECT -0.130 -0.075 0.420 0.075 ;
END VIA5_2CUT_E

# Via 9 - double cut west
VIA VIA5_2CUT_W DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal5 ;
    RECT -0.420 -0.075  0.130 0.075 ;
  LAYER Via5 ;
    RECT -0.360 -0.070 -0.220 0.070 ;
    RECT -0.070 -0.070  0.070 0.070 ;
  LAYER Metal6 ;
    RECT -0.420 -0.075  0.130 0.075 ;
END VIA5_2CUT_W

# Via 10 - double cut north
VIA VIA5_2CUT_N DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal5 ;
    RECT -0.075 -0.130 0.075 0.420 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT -0.070  0.220 0.070 0.360 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.420 ;
END VIA5_2CUT_N

# Via 11 - double cut south
VIA VIA5_2CUT_S DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal5 ;
    RECT -0.075 -0.420 0.075  0.130 ;
  LAYER Via5 ;
    RECT -0.070 -0.360 0.070 -0.220 ;
    RECT -0.070 -0.070 0.070  0.070 ;
  LAYER Metal6 ;
    RECT -0.075 -0.420 0.075  0.130 ;
END VIA5_2CUT_S

# Via 12 - quad cut square
VIA VIA5_2X2CUT DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal5 ;
    RECT -0.275 -0.220  0.275  0.220 ;
  LAYER Via5 ;
    RECT  0.075  0.075  0.215  0.215 ;
    RECT -0.215  0.075 -0.075  0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT  0.075 -0.215  0.215 -0.075 ;
  LAYER Metal6 ;
    RECT -0.220 -0.275  0.220  0.275 ;
END VIA5_2X2CUT


# Via 1 - Pin access Metal4 or Metal5
VIA VIA6X DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal7 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA6X

# Via 2 - Pin access Metal4 or Metal5
VIA VIA6H DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal7 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA6H

# Via 3 - Pin access Metal4 or Metal5
VIA VIA6V DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.130 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal7 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA6V

# Via 4 - Pin access Metal4 or Metal5
VIA VIA6XR90 DEFAULT
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.130 -0.075 0.130 0.075 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal7 ;
    RECT -0.075 -0.130 0.075 0.130 ;
END VIA6XR90

## Via 5 - TOS via for 5 signal wire (no pin access)
#VIA VIA6TOS DEFAULT
#  TOPOFSTACKONLY
#  RESISTANCE 1.4 ;
#  LAYER Metal6 ;
#    RECT -0.135 -0.170 0.135 0.170 ;
#  LAYER Via6 ;
#    RECT -0.070 -0.070 0.070 0.070 ;
#  LAYER Metal7 ;
#    RECT -0.130 -0.075 0.130 0.075 ;
#END VIA6TOS

VIA VIA6TOS DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.075 -0.27 0.075 0.27 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER Metal7 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA6TOS

VIA VIA6TOS_S DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.075 -0.41 0.075 0.13 ;
  LAYER Via6 ;
    RECT -0.070 -0.07 0.070 0.07 ;
  LAYER Metal7 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA6TOS_S

VIA VIA6TOS_N DEFAULT TOPOFSTACKONLY
  RESISTANCE 1.4 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.41 ;
  LAYER Via6 ;
    RECT -0.070 -0.07 0.070 0.07 ;
  LAYER Metal7 ;
    RECT -0.130 -0.075 0.130 0.075 ;
END VIA6TOS_N

# Via 6 - double cut north
VIA VIA6_2CUT_N DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal6 ;
    RECT -0.075 -0.130 0.075 0.420 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT -0.070  0.220 0.070 0.360 ;
  LAYER Metal7 ;
    RECT -0.075 -0.130 0.075 0.420 ;
END VIA6_2CUT_N

# Via 7 - double cut south
VIA VIA6_2CUT_S DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal6 ;
    RECT -0.075 -0.420 0.075  0.130 ;
  LAYER Via6 ;
    RECT -0.070 -0.360 0.070 -0.220 ;
    RECT -0.070 -0.070 0.070  0.070 ;
  LAYER Metal7 ;
    RECT -0.075 -0.420 0.075  0.130 ;
END VIA6_2CUT_S

# Via 8 - double cut east
VIA VIA6_2CUT_E DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal6 ;
    RECT -0.130 -0.075 0.420 0.075 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    RECT  0.220 -0.070 0.360 0.070 ;
  LAYER Metal7 ;
    RECT -0.130 -0.075 0.420 0.075 ;
END VIA6_2CUT_E

# Via 9 - double cut west
VIA VIA6_2CUT_W DEFAULT
  RESISTANCE 0.7 ;
  LAYER Metal6 ;
    RECT -0.420 -0.075  0.130 0.075 ;
  LAYER Via6 ;
    RECT -0.360 -0.070 -0.220 0.070 ;
    RECT -0.070 -0.070  0.070 0.070 ;
  LAYER Metal7 ;
    RECT -0.420 -0.075  0.130 0.075 ;
END VIA6_2CUT_W

# Via 10 - quad cut square
VIA VIA6_2X2CUT DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal6 ;
    RECT -0.220 -0.275  0.220  0.275 ;
  LAYER Via6 ;
    RECT  0.075  0.075  0.215  0.215 ;
    RECT -0.215  0.075 -0.075  0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT  0.075 -0.215  0.215 -0.075 ;
  LAYER Metal7 ;
    RECT -0.275 -0.220  0.275  0.220 ;
END VIA6_2X2CUT


# Via 1 - pin access via
VIA VIA7X DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal7 ;
    RECT -0.260 -0.210 0.260 0.210 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal8 ;
    RECT -0.230 -0.280 0.230 0.280 ;
END VIA7X

# Via 2 - pin access via
VIA VIA7V DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal7 ;
    RECT -0.210 -0.260 0.210 0.260 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal8 ;
    RECT -0.230 -0.280 0.230 0.280 ;
END VIA7V


# Via 3 - pin access via
VIA VIA7H DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal7 ;
    RECT -0.260 -0.210 0.260 0.210 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal8 ;
    RECT -0.280 -0.230 0.280 0.230 ;
END VIA7H

# Via 4 - pin access via
VIA VIA7XR90 DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal7 ;
    RECT -0.210 -0.260 0.210 0.260 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal8 ;
    RECT -0.230 -0.280 0.230 0.280 ;
END VIA7XR90

# Note, there are no VIA7TOS* vias because Metal7 already meets MAR rules.

# Via 5 - double cut east
VIA VIA7_2CUT_E DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal7 ;
    RECT -0.260 -0.210 0.980 0.210 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    RECT  0.540 -0.180 0.900 0.180 ;
  LAYER Metal8 ;
    RECT -0.280 -0.230 1.000 0.230 ;
END VIA7_2CUT_E

# Via 6 - double cut west
VIA VIA7_2CUT_W DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal7 ;
    RECT -0.980 -0.210  0.260 0.210 ;
  LAYER Via7 ;
    RECT -0.900 -0.180 -0.540 0.180 ;
    RECT -0.180 -0.180  0.180 0.180 ;
  LAYER Metal8 ;
    RECT -1.000 -0.230  0.280 0.230 ;
END VIA7_2CUT_W

# Via 7 - double cut north
VIA VIA7_2CUT_N DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal7 ;
    RECT -0.210 -0.260 0.210 0.980 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    RECT -0.180  0.540 0.180 0.900 ;
  LAYER Metal8 ;
    RECT -0.230 -0.280 0.230 1.000 ;
END VIA7_2CUT_N

# Via 8 - double cut south
VIA VIA7_2CUT_S DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal7 ; 
    RECT -0.210 -0.980 0.210  0.260 ;
  LAYER Via7 ;
    RECT -0.180 -0.900 0.180 -0.540 ;
    RECT -0.180 -0.180 0.180  0.180 ;
  LAYER Metal8 ;
    RECT -0.230 -1.000 0.230  0.280 ;
END VIA7_2CUT_S

# Via 9 - quad cut square
VIA VIA7_2X2CUT DEFAULT
  RESISTANCE 0.0875 ;
  LAYER Metal7 ;
    RECT -0.710 -0.660  0.710  0.660 ;
  LAYER Via7 ;
    RECT  0.270  0.270  0.630  0.630 ;
    RECT -0.630  0.270 -0.270  0.630 ;
    RECT -0.630 -0.630 -0.270 -0.270 ;
    RECT  0.270 -0.630  0.630 -0.270 ;
  LAYER Metal8 ;
    RECT -0.680 -0.730  0.680  0.730 ;
END VIA7_2X2CUT

# Via 1 - Signal routing via
VIA VIA8X DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal8 ;
    RECT -0.230 -0.260 0.230 0.260 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal9 ;
    RECT -0.280 -0.230 0.280 0.230 ;
END VIA8X

# Via 2 - Signal routing via
VIA VIA8H DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal8 ;
    RECT -0.260 -0.230 0.260 0.230 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal9 ;
    RECT -0.280 -0.230 0.280 0.230 ;
END VIA8H

# Via 3
VIA VIA8V DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal8 ;
    RECT -0.230 -0.260 0.230 0.260 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal9 ;
    RECT -0.230 -0.280 0.230 0.280 ;
END VIA8V

# Via 4 - Signal routing via
VIA VIA8XR90 DEFAULT
  RESISTANCE 0.35 ;
  LAYER Metal8 ;
    RECT -0.260 -0.230 0.260 0.230 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER Metal9 ;
    RECT -0.230 -0.280 0.230 0.280 ;
END VIA8XR90


# Via 8 - double cut east
VIA VIA8_2CUT_E DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal8 ;
    RECT -0.260 -0.230 0.980 0.230 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    RECT  0.540 -0.180 0.900 0.180 ;
  LAYER Metal9 ;
    RECT -0.280 -0.230 1.000 0.230 ;
END VIA8_2CUT_E

# Via 9 - double cut west
VIA VIA8_2CUT_W DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal8 ;
    RECT -0.980 -0.230  0.260 0.230 ;
  LAYER Via8 ;
    RECT -0.900 -0.180 -0.540 0.180 ;
    RECT -0.180 -0.180  0.180 0.180 ;
  LAYER Metal9 ;
    RECT -1.000 -0.230  0.280 0.230 ;
END VIA8_2CUT_W

# Via 10 - double cut north
VIA VIA8_2CUT_N DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal8 ;
    RECT -0.230 -0.260 0.230 0.980 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    RECT -0.180  0.540 0.180 0.900 ;
  LAYER Metal9 ;
    RECT -0.230 -0.280 0.230 1.000 ;
END VIA8_2CUT_N

# Via 11 - double cut south
VIA VIA8_2CUT_S DEFAULT
  RESISTANCE 0.175 ;
  LAYER Metal8 ;
    RECT -0.230 -0.980 0.230  0.260 ;
  LAYER Via8 ;
    RECT -0.180 -0.900 0.180 -0.540 ;
    RECT -0.180 -0.180 0.180  0.180 ;
  LAYER Metal9 ;
    RECT -0.230 -1.000 0.230  0.280 ;
END VIA8_2CUT_S

# Via 12 - quad cut square
VIA VIA8_2X2CUT DEFAULT
  RESISTANCE 0.0875 ;
  LAYER Metal8 ;
    RECT -0.660 -0.710  0.660  0.710 ;
  LAYER Via8 ;
    RECT  0.270  0.270  0.630  0.630 ;
    RECT -0.630  0.270 -0.270  0.630 ;
    RECT -0.630 -0.630 -0.270 -0.270 ;
    RECT  0.270 -0.630  0.630 -0.270 ;
  LAYER Metal9 ;
    RECT -0.730 -0.680  0.730  0.680 ;
END VIA8_2X2CUT



# SPECIAL NET ROUTING VIAS
VIA VIA1_2CUT_H
  RESISTANCE 0.7 ;
  LAYER Metal1 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via1 ;
    RECT -0.215 -0.070 -0.075 0.070 ;
    RECT  0.075 -0.070  0.215 0.070 ;
  LAYER Metal2 ;
    RECT -0.275 -0.075 0.275 0.075 ;
END VIA1_2CUT_H

VIA VIA1_2CUT_V
  RESISTANCE 0.7 ;
  LAYER Metal1 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via1 ;
    RECT -0.070 -0.215  0.070 -0.075 ;
    RECT -0.070  0.075  0.070 0.215 ;
  LAYER Metal2 ;
    RECT -0.075 -0.275 0.075 0.275 ;
END VIA1_2CUT_V

# Enforce the use of double cut vias
# First layer (primary direction) cover widths less than 3 via cuts
# Second layer cover widths from via width to 3 via cuts

VIARULE VIARULE1_2CUT_H
  LAYER Metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA1_2CUT_H ;
END VIARULE1_2CUT_H
    
VIARULE VIARULE1_2CUT_V
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA1_2CUT_V ;
END VIARULE1_2CUT_V

VIARULE VIA1ARRAY GENERATE
  LAYER Metal1 ;
    #DIRECTION HORIZONTAL
    ENCLOSURE .06 .005 ; 
    WIDTH 0.12 TO 12.00 ;
  LAYER Metal2 ;
    #DIRECTION VERTICAL
    ENCLOSURE .005 .06 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Via1 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    SPACING .34 BY .34 ;
    RESISTANCE 1.4 ;
END VIA1ARRAY        


VIA VIA2_2CUT_H
  RESISTANCE 0.7 ;
  LAYER Metal2 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via2 ;
    RECT -0.215 -0.070 -0.075 0.070 ;
    RECT  0.075 -0.070  0.215 0.070 ;
  LAYER Metal3 ;
    RECT -0.275 -0.075 0.275 0.075 ;
END VIA2_2CUT_H


VIA VIA2_2CUT_V
  RESISTANCE 0.7 ;
  LAYER Metal2 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via2 ;
    RECT -0.070 -0.215  0.070 -0.075 ;
    RECT -0.070  0.075  0.070 0.215 ;
  LAYER Metal3 ;
    RECT -0.075 -0.275 0.075 0.275 ;
END VIA2_2CUT_V

VIARULE VIARULE2_2CUT_H
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA2_2CUT_H ;
END VIARULE2_2CUT_H

VIARULE VIARULE2_2CUT_V
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA2_2CUT_V ;
END VIARULE2_2CUT_V


VIARULE VIA2ARRAY GENERATE
  LAYER Metal2 ;
    #DIRECTION VERTICAL ;
    ENCLOSURE .005 .06 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Metal3 ;
    #DIRECTION HORIZONTAL ;
    ENCLOSURE .06 .005 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Via2 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    SPACING .34 BY .34 ;
    RESISTANCE 1.4 ;
END VIA2ARRAY

VIA VIA3_2CUT_H
  RESISTANCE 0.7 ;
  LAYER Metal3 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via3 ;
    RECT -0.215 -0.070 -0.075 0.070 ;
    RECT  0.075 -0.070  0.215 0.070 ;
  LAYER Metal4 ;
    RECT -0.275 -0.075 0.275 0.075 ;
END VIA3_2CUT_H

VIA VIA3_2CUT_V
  RESISTANCE 0.7 ;
  LAYER Metal3 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via3 ;
    RECT -0.070 -0.215  0.070 -0.075 ;
    RECT -0.070  0.075  0.070 0.215 ;
  LAYER Metal4 ;
    RECT -0.075 -0.275 0.075 0.275 ;
END VIA3_2CUT_V

VIARULE VIARULE3_2CUT_H
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA3_2CUT_H ;
END VIARULE3_2CUT_H

VIARULE VIARULE3_2CUT_V
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA3_2CUT_V ;
END VIARULE3_2CUT_V


VIARULE VIA3ARRAY GENERATE
  LAYER Metal3 ;
    #DIRECTION HORIZONTAL ;
    ENCLOSURE .06 .005 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Metal4 ;
    #DIRECTION VERTICAL ;
    ENCLOSURE .005 .06 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Via3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    SPACING .34 BY .34 ;
    RESISTANCE 1.4 ;
END VIA3ARRAY

VIA VIA4_2CUT_H
  RESISTANCE 0.7 ;
  LAYER Metal4 ; 
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via4 ;
    RECT -0.215 -0.070 -0.075 0.070 ;
    RECT  0.075 -0.070  0.215 0.070 ;
  LAYER Metal5 ;
    RECT -0.275 -0.075 0.275 0.075 ;
END VIA4_2CUT_H

VIA VIA4_2CUT_V
  RESISTANCE 0.7 ;
  LAYER Metal4 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via4 ; 
    RECT -0.070 -0.215  0.070 -0.075 ;
    RECT -0.070  0.075  0.070 0.215 ;
  LAYER Metal5 ;
    RECT -0.075 -0.275 0.075 0.275 ;
END VIA4_2CUT_V

VIARULE VIARULE4_2CUT_H
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ; 
    WIDTH 0.55 TO 1.170 ;
  VIA VIA4_2CUT_H ;
END VIARULE4_2CUT_H

VIARULE VIARULE4_2CUT_V
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal5 ; 
    DIRECTION HORIZONTAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA4_2CUT_V ;
END VIARULE4_2CUT_V


VIARULE VIA4ARRAY GENERATE
  LAYER Metal4 ;
    #DIRECTION VERTICAL ;
    ENCLOSURE .005 .06 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Metal5 ;
    #DIRECTION HORIZONTAL ;
    ENCLOSURE .06 .005 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Via4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    SPACING .34 BY .34 ;
    RESISTANCE 1.4 ;
END VIA4ARRAY


VIA VIA5_2CUT_H
  RESISTANCE 0.7 ;
  LAYER Metal5 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via5 ;
    RECT -0.215 -0.070 -0.075 0.070 ;
    RECT  0.075 -0.070  0.215 0.070 ;
  LAYER Metal6 ;
    RECT -0.275 -0.075 0.275 0.075 ;
END VIA5_2CUT_H


VIA VIA5_2CUT_V
  RESISTANCE 0.7 ;
  LAYER Metal5 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via5 ;
    RECT -0.070 -0.215  0.070 -0.075 ;
    RECT -0.070  0.075  0.070 0.215 ;
  LAYER Metal6 ;
    RECT -0.075 -0.275 0.075 0.275 ;
END VIA5_2CUT_V

VIARULE VIARULE5_2CUT_H
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal6 ;
    DIRECTION VERTICAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA5_2CUT_H ;
END VIARULE5_2CUT_H

VIARULE VIARULE5_2CUT_V
  LAYER Metal6 ;
    DIRECTION VERTICAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA5_2CUT_V ;
END VIARULE5_2CUT_V


VIARULE VIA5ARRAY GENERATE
  LAYER Metal5 ;
    #DIRECTION HORIZONTAL
    ENCLOSURE .06 .005 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Metal6 ;
    #DIRECTION VERTICAL
    ENCLOSURE .005 .06 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Via5 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    SPACING .34 BY .34 ;
    RESISTANCE 1.4 ;
END VIA5ARRAY

VIA VIA6_2CUT_H
  RESISTANCE 0.7 ;
  LAYER Metal6 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via6 ;
    RECT -0.215 -0.070 -0.075 0.070 ;
    RECT  0.075 -0.070  0.215 0.070 ;
  LAYER Metal7 ;
    RECT -0.275 -0.075 0.275 0.075 ;
END VIA6_2CUT_H

VIA VIA6_2CUT_V
  RESISTANCE 0.7 ;
  LAYER Metal6 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via6 ;
    RECT -0.070 -0.215  0.070 -0.075 ;
    RECT -0.070  0.075  0.070 0.215 ;
  LAYER Metal7 ;
    RECT -0.075 -0.275 0.075 0.275 ;
END VIA6_2CUT_V

VIARULE VIARULE6_2CUT_H
  LAYER Metal7 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal6 ;
    DIRECTION VERTICAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA6_2CUT_H ;
END VIARULE6_2CUT_H

VIARULE VIARULE6_2CUT_V
  LAYER Metal6 ;
    DIRECTION VERTICAL ;
    WIDTH 0.12 TO 1.170 ;
  LAYER Metal7 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.55 TO 1.170 ;
  VIA VIA6_2CUT_V ;
END VIARULE6_2CUT_V


VIARULE VIA6ARRAY GENERATE
  LAYER Metal6 ;
    #DIRECTION VERTICAL ;
    ENCLOSURE .005 .06 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Metal7 ;
    #DIRECTION HORIZONTAL ;
    ENCLOSURE .06 .005 ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Via6 ;
    RECT -0.070 -0.070 0.070 0.070 ;
    SPACING .34 BY .34 ;
    RESISTANCE 1.4 ;
END VIA6ARRAY


VIA VIA7_2CUT_H
  RESISTANCE 0.175 ;
  LAYER Metal7 ;
    RECT -0.620 -0.210 0.620 0.210 ;
  LAYER Via7 ;
    RECT -0.540 -0.180 -0.180 0.180 ;
    RECT  0.180 -0.180  0.540 0.180 ;
  LAYER Metal8 ;
    RECT -0.640 -0.230 0.640 0.230 ;
END VIA7_2CUT_H
  
VIA VIA7_2CUT_V
  RESISTANCE 0.175 ;
  LAYER Metal7 ;
    RECT -0.210 -0.620 0.210 0.620 ;
  LAYER Via7 ;
    RECT -0.180 -0.540  0.180 -0.180 ;
    RECT -0.180  0.180  0.180  0.540 ;
  LAYER Metal8 ;
    RECT -0.230 -0.640 0.230 0.640 ;
END VIA7_2CUT_V
    
VIARULE VIARULE7_2CUT_H
  LAYER Metal7 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.14 TO 3.065 ;
  LAYER Metal8 ;
    DIRECTION VERTICAL ;
    WIDTH 1.28 TO 3.185 ;
  VIA VIA7_2CUT_H ;
END VIARULE7_2CUT_H
    
VIARULE VIARULE7_2CUT_V
  LAYER Metal8 ;
    DIRECTION VERTICAL ; 
    WIDTH 0.44 TO 3.065 ;
  LAYER Metal7 ;
    DIRECTION HORIZONTAL ;
    WIDTH 1.28 TO 3.185 ;
  VIA VIA7_2CUT_V ;
END VIARULE7_2CUT_V


VIARULE VIA7ARRAY GENERATE
  LAYER Metal7 ;
    #DIRECTION HORIZONTAL ;
    ENCLOSURE .08 .03  ;
    WIDTH 0.14 TO 12.00 ;
  LAYER Metal8 ;
    #DIRECTION VERTICAL ;
    ENCLOSURE .05 .10 ;
    WIDTH 0.44 TO 12.00 ;
  LAYER Via7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    SPACING .90 BY .90 ;    
    RESISTANCE 0.35 ;
END VIA7ARRAY

VIA VIA8_2CUT_H
  RESISTANCE 0.175 ;
  LAYER Metal8 ;
    RECT -0.620 -0.230 0.620 0.230 ;
  LAYER Via8 ;
    RECT -0.540 -0.180 -0.180 0.180 ;
    RECT  0.180 -0.180  0.540 0.180 ;
  LAYER Metal9 ;
    RECT -0.640 -0.230 0.640 0.230 ;
END VIA8_2CUT_H
  
VIA VIA8_2CUT_V
  RESISTANCE 0.175 ;
  LAYER Metal8 ;
    RECT -0.230 -0.620 0.230 0.620 ;
  LAYER Via8 ;
    RECT -0.180 -0.540  0.180 -0.180 ;
    RECT -0.180  0.180  0.180  0.540 ;
  LAYER Metal9 ;
    RECT -0.230 -0.640 0.230 0.640 ;
END VIA8_2CUT_V
    
VIARULE VIARULE8_2CUT_H
  LAYER Metal8 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.44 TO 3.065 ;
  LAYER Metal9 ;
    DIRECTION VERTICAL ;
    WIDTH 1.28 TO 3.185 ;
  VIA VIA8_2CUT_H ;
END VIARULE8_2CUT_H
    
VIARULE VIARULE8_2CUT_V
  LAYER Metal8 ;
    DIRECTION VERTICAL ; 
    WIDTH 0.44 TO 3.065 ;
  LAYER Metal9 ;
    DIRECTION HORIZONTAL ;
    WIDTH 1.28 TO 3.185 ;
  VIA VIA8_2CUT_V ;
END VIARULE8_2CUT_V

VIARULE VIA8ARRAY GENERATE
  LAYER Metal8 ;
    #DIRECTION VERTICAL ;
    ENCLOSURE .04 .08  ;
    #ENCLOSURE .03 .08  ; # .03 does not meet minimum Metal8 width
    WIDTH 0.44 TO 12.00 ;
  LAYER Metal9 ;
    #DIRECTION HORIZONTAL ;
    ENCLOSURE .10 .05  ;
    WIDTH 0.44 TO 12.00 ;
  LAYER Via8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
    SPACING .90 BY .90 ;    
    RESISTANCE 0.35 ;
END VIA8ARRAY           
#
#
#
#MACRO statement...
#   PIN statement...
#   OBS statement...

#BEGINEXT "tag-in-quotes"
#   extension statements
#ENDEXT

END LIBRARY
